��,�      }�(�database��editorCode.database��Database���)��}�(�bodies�]��$editorCode.shapeInternals.editorBody��
BodyStatic���)��}�(�label��Level��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G@WP��b�h!G@JM��)ubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@Y�v'��h!G@O�x�R��ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G@f汆3��r0c1�G�       �r0c2�G@W4fwOh�r1c0�G        �r1c1�G@f汆3��r1c2�G@I����B�ub�objectAnchor�h)��}�(h G@W4fwOhh!G@I����B�ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G@f汆3�ub�shapes�]�(�%editorCode.shapeInternals.editorShape��Line���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@2�3��YTh!G?���5�ٰububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@;V��x�Lh!G@$�It��ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��type��Line��internal��)editorCode.shapeInternals.editorShapeSpec��LineSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G�.��+?ڸh!G�":�f$pTubh"h)��}�(h G� ������h!G�"�u	(ububh)��}�(hh)��}�(h G�)5��9��h!G�"M��g�ubh"h)��}�(h G@"��@�}h!G�"}6��ububh)��}�(hh)��}�(h G�%��V�-h!G�!�hYp<�ubh"h)��}�(h G@4XAM��h!G����5��ububh)��}�(hh)��}�(h G�$U�_��Fh!G�!6h��ubh"h)��}�(h G@9_����h!G��FDA�Pububh)��}�(hh)��}�(h G�#+ж>h!G� ��r��ubh"h)��}�(h G@=h*�J��h!G��d�J��ububh)��}�(hh)��}�(h G�"u�?�Ih!G� `�ȶ�rubh"h)��}�(h G@?�
!�h!G�--�
R@ububh)��}�(hh)��}�(h G�!+g�WKh!G���r���ubh"h)��}�(h G@A�s����h!G?܋!�q� ububh)��}�(hh)��}�(h G� K��w�h!G�m��=�&ubh"h)��}�(h G@CZ=�/Ԟh!G@�
�uIPububh)��}�(hh)��}�(h G�����Yh!G�M�#ubh"h)��}�(h G@D:�>s��h!G@�Pr�K�ububh)��}�(hh)��}�(h G���Y�H�h!G��v��ubh"h)��}�(h G@E��y�~h!G@!/ܠ��ububh)��}�(hh)��}�(h G�=(C&h!G��c���ubh"h)��}�(h G@Gr�~�h!G@&�[6,(ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��LinePhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G�%��H)oh!G� �ԔHub�user�h)��}�(h G        h!G        ubh"h)��}�(h G�%��H)oh!G� �ԔHub�userDefined��ub�area�G?�PsBBG�density�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      hˉub�mass�h�)��}�(h�G?�      h�G        h"G?�PsBBG�hˉub�moment�h�)��}�(h�G?�����'�h�G        h"G?�����'�hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@Rn,�rh!G?��z+u��ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@>�"��{h!G@"��!�Jubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1�hfhghhhk)��}�(hn]�(h)��}�(hh)��}�(h G�~ 8�*h!G�>Sp��ubh"h)��}�(h G@G	��m0h!G@&Ln�p�ububh)��}�(hh)��}�(h G�	,�$2�h!G�f��H/�ubh"h)��}�(h G@FI���śh!G@Y3 &�ububh)��}�(hh)��}�(h G�����h!G�Ԭյ�bubh"h)��}�(h G@E���ӷh!G@�NR�8ububh)��}�(hh)��}�(h G�䚑���h!G����7�ubh"h)��}�(h G@E�����h!G?� ��g ububh)��}�(hh)��}�(h G��H�Sh!G� /j� �ubh"h)��}�(h G@F��h!G�V�@ ububh)��}�(hh)��}�(h G��}\�zh!G�!�G���ubh"h)��}�(h G@L;�A�?Eh!G�6e��ububh)��}�(hh)��}�(h G���ׇ-�h!G�!��t��!ubh"h)��}�(h G@O�)���h!G���PP�ububh)��}�(hh)��}�(h G�Cn
J�h!G� �����ubh"h)��}�(h G@R�^�\",h!G���22��ububh)��}�(hh)��}�(h G?�iH|Z�h!G�!(}�v�ubh"h)��}�(h G@X�*�h!G��O��@ububh)��}�(hh)��}�(h G?�}���ph!G� U��zX�ubh"h)��}�(h G@Y��[���h!G�	�j6րububh)��}�(hh)��}�(h G?�� �\8h!G��&V�p�ubh"h)��}�(h G@Z����h!G?�Λ%܀ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G��s��s�h!G� �ғ��ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��s��s�h!G� �ғ��ubhˉubh�G?ΰ�_�h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?ΰ�_�hˉubh�h�)��}�(h�G@�AI�h�G        h"G@�AI�hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@b�.�3�Fh!G@?rd��ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@G1T~ggh!G@/���ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfhghhhk)��}�(hn]�(h)��}�(hh)��}�(h G?��/aԈh!G����GQ{ubh"h)��}�(h G@Z��[�h!G?�`��0�ububh)��}�(hh)��}�(h G?�m�>)i�h!G�"��&�a�ubh"h)��}�(h G@Z(0��qh!G�$<Lׇ�@ububh)��}�(hh)��}�(h G@��P2h!G�"�"�:ubh"h)��}�(h G@[&"%Wh!G�$�͔.��ububh)��}�(hh)��}�(h G@�m:']h!G�"���+8ubh"h)��}�(h G@_S�#�h!G�$�䢁CLububh)��}�(hh)��}�(h G@���h!G�"�D*��ubh"h)��}�(h G@aÙjFيh!G�$��M ububh)��}�(hh)��}�(h G@&��]Ƌ�h!G�"�fdBrubh"h)��}�(h G@d�V��hh!G�%�s��|ububh)��}�(hh)��}�(h G@)x�h!G�"M5�^3.ubh"h)��}�(h G@fV�"Eh!G�"}ۓ
�Dububh)��}�(hh)��}�(h G@*��|+�h!G�!tp��Xubh"h)��}�(h G@f��:��,h!G��&��G�ububh)��}�(hh)��}�(h G@,\3���h!G� �Y�:6ubh"h)��}�(h G@gB�]��h!G�����2t�ububh)��}�(hh)��}�(h G@- S��9h!G��*m
�ubh"h)��}�(h G@g�]Dߐ,h!G?���x� ububh)��}�(hh)��}�(h G@.z�m;^h!G��">J�wubh"h)��}�(h G@h"6�1sh!G@�h�2�Hububh)��}�(hh)��}�(h G@/� ���dh!G�����ubh"h)��}�(h G@h���� h!G@4M٫���ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G@"2����gh!G�!'�`ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@"2����gh!G�!'�`ubhˉubh�G?ׅb���h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?ׅb���hˉubh�h�)��}�(h�G@!��Q�
h�G        h"G@!��Q�
hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@WO���kh!G@Q���Sububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@Y��,Ue<h!G@G�]�&Jubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hf�Line�hhhk)��}�(hn]�(h)��}�(hh)��}�(h G@/��C��<h!G��l|`טubh"h)��}�(h G@h�����h!G@4 �����ububh)��}�(hh)��}�(h G@/��ܹ2�h!G@jܝ�ġubh"h)��}�(h G@h�}f�dsh!G@SD��\+ububh)��}�(hh)��}�(h G@,����h!G@����zubh"h)��}�(h G@gq*���h!G@WP��F@ububh)��}�(hh)��}�(h G@(�.(��
h!G@�'Pҫ�ubh"h)��}�(h G@e��dph!G@Y�`��?ububh)��}�(hh)��}�(h G@)Pk�2h!G@"7k��A�ubh"h)��}�(h G@a�=�#��h!G@[�v�b�ububh)��}�(hh)��}�(h G@�M�`��h!G@"�Yޘ�ubh"h)��}�(h G@]�Hށlh!G@\e�c�O ububh)��}�(hh)��}�(h G?�Ծ��_h!G@#���-ubh"h)��}�(h G@Y*�W�ʿh!G@\�����xububh)��}�(hh)��}�(h G�-Y���h!G@#aG*l�pubh"h)��}�(h G���c�ϰh!G@\�5����ububh)��}�(hh)��}�(h G�.�講>h!G@"�C��b�ubh"h)��}�(h G�!����Xh!G@\_>.���ububh)��}�(hh)��}�(h G�/9v�J�h!G@!y�M��kubh"h)��}�(h G�%!Ulֈh!G@[4�ݾnububh)��}�(hh)��}�(h G�/%ewʋ�h!G@�L0:G<ubh"h)��}�(h G�$��>��h!G@X�F�4ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G@�bC���h!G@Ro>�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@�bC���h!G@Ro>�ubhˉubh�G?�n��t��h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�n��t��hˉubh�h�)��}�(h�G@^�8V�ah�G        h"G@^�8V�ahˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G�
v�MQ�ph!G@S�t��ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@<�՝�h!G@4 ��5�Aubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_4�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G�/$�+'M�h!G@�O�R|ubh"h)��}�(h G�$�d����h!G@X���kE�ububh)��}�(hh)��}�(h G�.��(�1h!G@��P��ubh"h)��}�(h G�"_^���xh!G@W��� ��ububh)��}�(hh)��}�(h G�-Ԇ����h!G@
`m��ubh"h)��}�(h G��\<���h!G@W�u�6�ububh)��}�(hh)��}�(h G�,x.�7��h!G@���vZ�ubh"h)��}�(h G��}�#� h!G@V�����ububh)��}�(hh)��}�(h G�*�F��ah!G@�U�G��ubh"h)��}�(h G@�]�`h!G@V+U�@�ububh)��}�(hh)��}�(h G�/*v	�~�h!G@PH_��ubh"h)��}�(h G�$�>"�h!G@U�X��ububh)��}�(hh)��}�(h G�/��H��h!G?��tk5<ubh"h)��}�(h G�$9��.W�h!G@M4�٠�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G�.�˖�Jh!G@�U'�^ubh�h)��}�(h G        h!G        ubh"h)��}�(h G�.�˖�Jh!G@�U'�^ubhˉubh�G?�<�,CVh�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�<�,CVhˉubh�h�)��}�(h�G?ⰾKI��h�G        h"G?ⰾKI��hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@A����=h!G@8�Wj|�ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@F��ɡ|�h!G@@��T�n�ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_5�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G�/�����h!G?� }�'�ubh"h)��}�(h G�$���pHh!G@M	�o�ububh)��}�(hh)��}�(h G�+v�ԏZh!G?��ab{�ubh"h)��}�(h G?�� �='�h!G@Kc�ׂububh)��}�(hh)��}�(h G�)vYR	!h!G?��a�G7�ubh"h)��}�(h G@ ��'3�h!G@I�`-Oqububh)��}�(hh)��}�(h G�#��*�h!G��]��	�0ubh"h)��}�(h G@=�D��.h!G@Fۏ��O�ububh)��}�(hh)��}�(h G��Z݁8
h!G��ԂC�ubh"h)��}�(h G@Kx�ҏ�h!G@E���J�ububh)��}�(hh)��}�(h G����1�Lh!G��JbO<ubh"h)��}�(h G@L8�mh!G@E��{�@ububh)��}�(hh)��}�(h G����2b��h!G��%�s�vPubh"h)��}�(h G@T&���%mh!G@H-ReC~�ububh)��}�(hh)��}�(h G�	|�P�h!G��:]΂oLubh"h)��}�(h G@P���3v�h!G@F $p�iububh)��}�(hh)��}�(h G��e�9�h!G���.��Wubh"h)��}�(h G@K�`�G�|h!G@D�pw�1�ububh)��}�(hh)��}�(h G�mDŵ�-h!G��K��w%�ubh"h)��}�(h G@J�K���h!G@Dţ_�uububh)��}�(hh)��}�(h G�"��S��6h!G��4����zubh"h)��}�(h G@?Dþ��h!G@D�M�\��ububh)��}�(hh)��}�(h G�(N��OUh!G���~`fubh"h)��}�(h G@(�FYU�Ph!G@F^a+ububh)��}�(hh)��}�(h G�/)?gˆ�h!G?�CI�=n@ubh"h)��}�(h G�$��{�hh!G@J��ֿl�ububh)��}�(hh)��}�(h G�/)�gc\h!G�!�zd7�ubh"h)��}�(h G�$��"��h!G���Xr`ububh)��}�(hh)��}�(h G�.�qY	D/h!G�"D�7�ubh"h)��}�(h G�!뾼
�h!G�"F�}��\ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G�$ꩥ�V�h!G��L����hubh�h)��}�(h G        h!G        ubh"h)��}�(h G�$ꩥ�V�h!G��L����hubhˉubh�G?�h� ��h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�h� ��hˉubh�h�)��}�(h�G@3��y��h�G        h"G@3��y��hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@V
Bhw-�h!G@)���Vpububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@дkɬ�h!G@�;�kpubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_6�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G���ĎM�h!G�I=UX]\ubh"h)��}�(h G@T=7!���h!G@�e�
��ububh)��}�(hh)��}�(h G?��Ej�/Ph!G�N�K&t[ubh"h)��}�(h G@W�M�3�mh!G@V�=�Apububh)��}�(hh)��}�(h G��J��Bm�h!G���b���ubh"h)��}�(h G@U� "Uamh!G@ �A�^Fububh)��}�(hh)��}�(h G���n�U��h!G�C�_�F\ubh"h)��}�(h G@T?���$h!G@���m�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G��y�_��h!G�^S�{ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��y�_��h!G�^S�{ubhˉubh�G?�t��>T�h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�t��>T�hˉubh�h�)��}�(h�G?�U��Oc�h�G        h"G?�U��Oc�hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@aC:!v�h!G@1N_�P(ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@=���/4h!G@,��h���ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_7�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G@Q���$h!G����6�ubh"h)��}�(h G@[Lmanh!G@%P��ôububh)��}�(hh)��}�(h G@	�QC�y�h!G�˺u��ubh"h)��}�(h G@\mR#�tnh!G@
��zspububh)��}�(hh)��}�(h G@&�����Hh!G�^�t��vubh"h)��}�(h G@d�����h!G@��Z�=�ububh)��}�(hh)��}�(h G@&����4h!G�����<ubh"h)��}�(h G@d����<�h!G@?�Ó��ububh)��}�(hh)��}�(h G@#���`�h!G���!�Pubh"h)��}�(h G@cɞ�:�h!G@7�Ls���ububh)��}�(hh)��}�(h G@�� �ueh!G��3O;�ubh"h)��}�(h G@a���uDh!G@2SDO���ububh)��}�(hh)��}�(h G@�y�*6h!G��G���ubh"h)��}�(h G@_����h!G@+t��#�@ububh)��}�(hh)��}�(h G@�"Յ��h!G���BG�_ubh"h)��}�(h G@[0����"h!G@%V�:�z�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G@��O�=�h!G���s�X�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@��O�=�h!G���s�X�ubhˉubh�G?�I2)R%h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�I2)R%hˉubh�h�)��}�(h�G@C7��`�h�G        h"G@C7��`�hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@g+zSsn2h!G@@I
dububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��x4��h!G@'��v���ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_8�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G@,��$�Ѫh!G�m��'subh"h)��}�(h G@g[ICۣ�h!G@4����Tububh)��}�(hh)��}�(h G@,���F�,h!G��a;�Tubh"h)��}�(h G@gV����2h!G@F2��'D�ububh)��}�(hh)��}�(h G@+�;��:h!G���l�`�ubh"h)��}�(h G@f��c8�h!G@>��u�(ububh)��}�(hh)��}�(h G@,���F�,h!G� ;�.��ubh"h)��}�(h G@gV����2h!G@5>uU���ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G@,X��Nh!G�iw�4��ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@,X��Nh!G�iw�4��ubhˉubh�G?�ㅄ�h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�ㅄ�hˉubh�h�)��}�(h�G?�7/���h�G        h"G?�7/���hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@fs�w�~h!G@G8�>U4tububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@~Z�h!G@����dubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_9�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G@),`�^�h!G��l���3ubh"h)��}�(h G@e�;�( .h!G@F��1p�ububh)��}�(hh)��}�(h G@+؂�6�h!G?�x7tl�hubh"h)��}�(h G@gT�j�.h!G@J� 2Q��ububh)��}�(hh)��}�(h G@(�fURjzh!G��6c�qqubh"h)��}�(h G@e�<��h!G@C��JX�hububh)��}�(hh)��}�(h G@)]��\h!G����o4�ubh"h)��}�(h G@e�ɘ��Fh!G@F�� 0��ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G@*/ v���h!G�������ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@*/ v���h!G�������ubhˉubh�G?����h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?����hˉubh�h�)��}�(h�G?�k�fZ��h�G        h"G?�k�fZ��hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@6������h!G@Tk�D��ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@��6'�h!G@�'��ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_10�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G�$�k��.lh!G@��ojU�ubh"h)��}�(h G@7K���Lh!G@V%����tububh)��}�(hh)��}�(h G�&#��R"<h!G@��c�a@ubh"h)��}�(h G@3k���Xh!G@Vwl�ububh)��}�(hh)��}�(h G�&��z;�h!G@��g_݊ubh"h)��}�(h G@0��ʦLh!G@U��Ti��ububh)��}�(hh)��}�(h G�'{����h!G@�H���ubh"h)��}�(h G@-��2�. h!G@T�¦Ttububh)��}�(hh)��}�(h G�'b¨c`h!G@��$z�ubh"h)��}�(h G@.���48h!G@S����ububh)��}�(hh)��}�(h G�&3H���h!G@)�K�;�ubh"h)��}�(h G@38��пph!G@R�Ş���ububh)��}�(hh)��}�(h G�$xt���h!G@�w�{�ubh"h)��}�(h G@8�����h!G@R���?�ububh)��}�(hh)��}�(h G�#XvE�h!G@��흚ubh"h)��}�(h G@<�{yXh!G@SO��7ububh)��}�(hh)��}�(h G�"߰̐�rh!G@+��x�ubh"h)��}�(h G@>3��(4h!G@S�'PYʽububh)��}�(hh)��}�(h G�"��o2�h!G@'i����ubh"h)��}�(h G@>z��_*�h!G@T��5�R�ububh)��}�(hh)��}�(h G�#�D.�F,h!G@�~�Q��ubh"h)��}�(h G@;|!�Lh!G@U�'��ububh)��}�(hh)��}�(h G�$ی��nh!G@��c�a@ubh"h)��}�(h G@7���}�h!G@Vwl�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G�%+���	Uh!G@o�M��ubh�h)��}�(h G        h!G        ubh"h)��}�(h G�%+���	Uh!G@o�M��ubhˉubh�G?H]r;�h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?H]r;�hˉubh�h�)��}�(h�G?�6�6{�h�G        h"G?�6�6{�hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@D#ɩ2h!G@U�	�^]�ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@
Y�<�hh!G@l��Y0ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_11�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G��j�L�h!G@�0�'ubh"h)��}�(h G@D�iCWh!G@V�m��&ububh)��}�(hh)��}�(h G� �����h!G@�kT���ubh"h)��}�(h G@B���8�h!G@V9�#�ububh)��}�(hh)��}�(h G� �@V��"h!G@�
�y��ubh"h)��}�(h G@B~7˔4|h!G@Uۗ���ububh)��}�(hh)��}�(h G� ��?`�Bh!G@���?�ubh"h)��}�(h G@B���7�h!G@UV���ububh)��}�(hh)��}�(h G�7)��]Qh!G@΢����ubh"h)��}�(h G@D}6-jG�h!G@T��&�ububh)��}�(hh)��}�(h G��+�)�h!G@���?�ubh"h)��}�(h G@E�'SWh!G@UV���ububh)��}�(hh)��}�(h G���Oz2h!G@����d$ubh"h)��}�(h G@E�[����h!G@V�Y��ububh)��}�(hh)��}�(h G��A��/h!G@��Ҽubh"h)��}�(h G@D+s�RD{h!G@V��T��ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G�����h!G@�E�`�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G�����h!G@�E�`�ubhˉubh�G?��283'h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?��283'hˉubh�h�)��}�(h�G?�Z  h�G        h"G?�Z  hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@Igtd(�<h!G@U�(��Kfububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@
1BR��(h!G@ i�\���ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_12�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G�>�1I�h!G@�N��ubh"h)��}�(h G@G�`>�#jh!G@V!QI�ububh)��}�(hh)��}�(h G��@G��h!G@�ݣ珊ubh"h)��}�(h G@I�Mh!G@UN�ͽ<�ububh)��}�(hh)��}�(h G�F2 9jLh!G@#z��Tubh"h)��}�(h G@K
��Sh!G@VUx3�Y�ububh)��}�(hh)��}�(h G�"��k�h!G@��~n�ubh"h)��}�(h G@Gں00�h!G@V*�`�kububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G�,�r�
h!G@:���9�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G�,�r�
h!G@:���9�ubhˉubh�G?��n�V�h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?��n�V�hˉubh�h�)��}�(h�G?x�݇aY�h�G        h"G?x�݇aY�hˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@PX
�N�@h!G@V��̟ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�*5P�h!G@k��8ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_13�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G�����h!G@�ߖ�l�ubh"h)��}�(h G@O��� h�h!G@Wp��qPububh)��}�(hh)��}�(h G�n%&B�$h!G@�I���ubh"h)��}�(h G@N6os���h!G@V�:c ��ububh)��}�(hh)��}�(h G���B��@h!G@� ���ubh"h)��}�(h G@M؏��8Fh!G@V:����ububh)��}�(hh)��}�(h G����_A�h!G@����}ubh"h)��}�(h G@N��wH�h!G@UbC቗zububh)��}�(hh)��}�(h G���{��h!G@��"�+ubh"h)��}�(h G@O��Q2h!G@T���l�ububh)��}�(hh)��}�(h G��P��Lh!G@)&�lubh"h)��}�(h G@Q'�y��uh!G@T���c�Rububh)��}�(hh)��}�(h G�	���h!G@�,˰�ubh"h)��}�(h G@Q��-��]h!G@UN&=�%
ububh)��}�(hh)��}�(h G�
!^�ʴ�h!G@�0��ubh"h)��}�(h G@Q�k~��Yh!G@V</���ububh)��}�(hh)��}�(h G���yo�h!G@d(�o��ubh"h)��}�(h G@P����/�h!G@V��y�Eububh)��}�(hh)��}�(h G���sw�qh!G@� ���ubh"h)��}�(h G@O�HQ�9�h!G@WwUPL� ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G��F���h!G@-�m�nxubh�h)��}�(h G        h!G        ubh"h)��}�(h G��F���h!G@-�m�nxubhˉubh�G?�h�m/�h�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G?�h�m/�hˉubh�h�)��}�(h�G?��C��jh�G        h"G?��C��jhˉubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@X��N��h!G@N��`�ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@U����+,h!G@A�\�Q�ubububh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G�       h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_14�hfj�  hhhk)��}�(hn]�(h)��}�(hh)��}�(h G@�ŎmB�h!G@pU:���ubh"h)��}�(h G@[���?�Dh!G@X��g�vububh)��}�(hh)��}�(h G��M�����h!G@�DW�ݪubh"h)��}�(h G@T�)��h!G@X5'�hjububh)��}�(hh)��}�(h G@���}(�h!G@�"��ubh"h)��}�(h G@\R���h!G@W$����ububh)��}�(hh)��}�(h G?j4��� h!G@� \T�$ubh"h)��}�(h G@W ��$�h!G@Ryw��x�ububh)��}�(hh)��}�(h G��,&�YLh!G?�s�J�,�ubh"h)��}�(h G@I�GNLSh!G@O=M
�Kububh)��}�(hh)��}�(h G�'l��<PLh!G?�z�ĵ_�ubh"h)��}�(h G@.\�a�.�h!G@O>ĊV��ububh)��}�(hh)��}�(h G�!`T�"�h!G?��}��ubh"h)��}�(h G@A�����h!G@N���ububh)��}�(hh)��}�(h G����=�Rh!G?�uu��/<ubh"h)��}�(h G@DY>��h!G@N ����ububh)��}�(hh)��}�(h G�#��߱@h!G?��4��ubh"h)��}�(h G@K&�x^h!G@N4c�/^ububh)��}�(hh)��}�(h G���)`h!G?��L���&ubh"h)��}�(h G@Ql�TToh!G@N����5ububh)��}�(hh)��}�(h G?��U�V��h!G@�ͻ��eubh"h)��}�(h G@W��!�Qh!G@Q��+ۛububh)��}�(hh)��}�(h G?�^w$�C�h!G@xq?t�ubh"h)��}�(h G@Z[hhE�h!G@S�I�̮�ububh)��}�(hh)��}�(h G@>��x�h!G@�B��lubh"h)��}�(h G@]'n
�5�h!G@V�@�=�:ububh)��}�(hh)��}�(h G@>_�G�~h!G@8�ir�ubh"h)��}�(h G@a̕�p�<h!G@U!%-Y�ububh)��}�(hh)��}�(h G@"� m�ԋh!G@�Tn�ubh"h)��}�(h G@c3ҵ[�>h!G@T����ububh)��}�(hh)��}�(h G@Q�Ր@�h!G?���f�vubh"h)��}�(h G@af�	h!G@MG���@ububh)��}�(hh)��}�(h G@N�ϩ�h!G��@�C@�ubh"h)��}�(h G@\��gc��h!G@E�,O��ububh)��}�(hh)��}�(h G����炉8h!G���A�ubh"h)��}�(h G@T��D��h!G@A��h��ububh)��}�(hh)��}�(h G� ����Oh!G�
���&��ubh"h)��}�(h G@B�R����h!G@=6�$u/lububh)��}�(hh)��}�(h G�(y���5h!G��.��ːubh"h)��}�(h G@'l�®�h!G@:s*�Z�ububh)��}�(hh)��}�(h G�uV!�h!G����@�rubh"h)��}�(h G@E{H��>h!G@:�e�<Z�ububh)��}�(hh)��}�(h G���^��h!G�	c��@��ubh"h)��}�(h G@Rp�V1�h!G@>4�88Q�ububh)��}�(hh)��}�(h G���Oj|*h!G���N�z_ubh"h)��}�(h G@T�н�h!G@?�]�|��ububh)��}�(hh)��}�(h G@�����h!G��Ý�� ubh"h)��}�(h G@^h�H�:�h!G@C^�َ-$ububh)��}�(hh)��}�(h G@���]5�h!G����7ف�ubh"h)��}�(h G@^��v���h!G@CB�f�ububh)��}�(hh)��}�(h G@�6�c`h!G?�5���ubh"h)��}�(h G@b$���h!G@KVj����ububh)��}�(hh)��}�(h G@&��ނ+h!G@J	!B�ubh"h)��}�(h G@e<�U��h!G@R�p�6Dububh)��}�(hh)��}�(h G@*g���9�h!G@����ubh"h)��}�(h G@ft"z��h!G@Q���݌Cububh)��}�(hh)��}�(h G@,Kr����h!G@���E�:ubh"h)��}�(h G@g;��Vh!G@PxG�2�ububh)��}�(hh)��}�(h G@,65���Nh!G@[IV[K�ubh"h)��}�(h G@g2�@�h!G@Q�,\}$ububh)��}�(hh)��}�(h G@*栁Gp�h!G@��[���ubh"h)��}�(h G@f�����h!G@R����=%ububh)��}�(hh)��}�(h G@(�%����h!G@kh��șubh"h)��}�(h G@e���n}�h!G@S�~�w��ububh)��}�(hh)��}�(h G@$����Ih!G@P�$ubh"h)��}�(h G@d7��^�)h!G@U�}4$�ububh)��}�(hh)��}�(h G@!>f��Egh!G@�u]� �ubh"h)��}�(h G@b���>#h!G@Uچ�owzububh)��}�(hh)��}�(h G@H�(��h!G@e;�ubh"h)��}�(h G@\!|m�`�h!G@X�rt�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G?�jH:���h!G?�^f���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?�jH:���h!G?�^f���ubhˉubh�G@^��Qmh�h�)��}�(h�G?�      h�G        h"G?�      hˉubh�h�)��}�(h�G?�      h�G        h"G@^��Qmhˉubh�h�)��}�(h�G@`ց�8�h�G        h"G@`ց�8�hˉubububehf�Static�h��+editorCode.shapeInternals.editorBodyPhysics��BodyStaticPhysics���)��}�(h�h�)��}�(h�h)��}�(h G        h!G        ubh�h)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubhˉubh�G?�      h�h�)��}�(h�G?�      h�G        h"G        hˉubh�h�)��}�(h�G?�      h�G        h"G        hˉubh�h�)��}�(h�G?�      h�G        h"G        hˉubububa�	shapeList�]�(hMh�jH  j�  j/  j�  j  jU  j�  j�  j?  j�  j  jY  j�  e�constraints�]��mappings�]��editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G@f汆3�h7G        h8G@W4fwOhh9G        h:G@f汆3�h;G@I����B�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�0      h!G�#�     ubh"h)��}�(h G�*=�Xw!�h!G�-~࢖�ububh)��}�(hh)��}�(h G@0      h!G�#�     ubh"h)��}�(h G@h�����h!G�-~࢖�ububh)��}�(hh)��}�(h G�0      h!G@#�     ubh"h)��}�(h G�*=�Xw!�h!G@]C��<  ububh)��}�(hh)��}�(h G@0      h!G@#�     ubh"h)��}�(h G@h�����h!G@]C��<  ubube�textureSize�]�(M Me�anchor�]�(G@�      G@s�     e�mappingSize�]�(M Me�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@�      h!G@s�     ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@W4fwOhh!G@I����B�ubububaub�textureSizes�]�(M M��K K ��j%  j%  j%  j%  j%  j%  j%  j%  j%  j%  j%  j%  j%  j%  e�texturePaths�]�(�data/textures/map02.png�� �j)  j)  j)  j)  j)  j)  j)  j)  j)  j)  j)  j)  j)  j)  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�h�currentShape�jH  �currentConstraint�N�currentMapping�j�  �currentMappingChannel�K hh)��}�(hhj�  j�  j�  j�  j�  j�  ububhj@  �object�h�prevCurrent�Nubj0  �ComSetBodyAsCurrent���)��}�(j5  j9  h�BODY��prev�hubj0  �ComRenameBody���)��}�(j�  hhj@  �newName�h�oldName�jH  ubj0  �ComLoadTexture���)��}�(hj@  �newPath�j(  �destChannel�K �newSize�j$  �oldPath�j)  �oldSize�j%  ubj0  �ComAddNewShape���)��}�(j5  j9  hj@  �shape�hM�	prevShape�Nj�  hubj0  �ComNewShapeAddPoint���)��}�(j]  hM�point�hpubj`  )��}�(j]  hMjc  hvubj`  )��}�(j]  hMjc  h|ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubj`  )��}�(j]  hMjc  h�ubjZ  )��}�(j5  j9  hj@  j]  h�j^  hMj�  hubj`  )��}�(j]  h�jc  h�ubj`  )��}�(j]  h�jc  h�ubj`  )��}�(j]  h�jc  j   ubj`  )��}�(j]  h�jc  j  ubj`  )��}�(j]  h�jc  j  ubj`  )��}�(j]  h�jc  j  ubj`  )��}�(j]  h�jc  j  ubj`  )��}�(j]  h�jc  j  ubj`  )��}�(j]  h�jc  j$  ubj`  )��}�(j]  h�jc  j*  ubj`  )��}�(j]  h�jc  j0  ubjZ  )��}�(j5  j9  hj@  j]  jH  j^  h�j�  hubj`  )��}�(j]  jH  jc  jd  ubj`  )��}�(j]  jH  jc  jj  ubj`  )��}�(j]  jH  jc  jp  ubj`  )��}�(j]  jH  jc  jv  ubj`  )��}�(j]  jH  jc  j|  ubj`  )��}�(j]  jH  jc  j�  ubj`  )��}�(j]  jH  jc  j�  ubj`  )��}�(j]  jH  jc  j�  ubj`  )��}�(j]  jH  jc  j�  ubj`  )��}�(j]  jH  jc  j�  ubj`  )��}�(j]  jH  jc  j�  ubj`  )��}�(j]  jH  jc  j�  ubj0  �ComStartTransform���)��}�(h,�editorCode.editorViewTransform��ContinuousTransform���)��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�
mouseParam��editorCode.editorMousePivot��MousePivotParams���)��}�(�pivot�h)��}�(h K h!K ub�begin�h)��}�(h G����`h!G��H�5l-@ub�end�h)��}�(h G��e�G���h!G���e� ub�dPivot�h)��}�(h G��e�G���h!G���e� ub�dEnd�h)��}�(h G��]�� h!G��iI}f ub�dA�hA)��}�(hDG?�[�Ev@hEG?�X�6@P�hFG?��%��ڦub�dS�G?�
`b�!�angleOffset�G� �#E�j��length�G?�ح���'ub�mode�K�active���obj�hub�newObj�h�
startPoint�h)��}�(h G����`h!G��H�5l-@ubj�  h)��}�(h K h!K ubj�  K�	processed���oldObjectAnchor�h)��}�(h G        h!G        ub�oldObjectAngle�hA)��}�(hDG        hEG        hFG?�      ub�oldObjectScale�G?�      ubj�  )��}�(h,j�  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G@, ���z\h!G@y�8K/�ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  j�  )��}�(j�  h)��}�(h G��t?�լ h!G?�U�ٺ� ubj�  h)��}�(h G@;�R#Nh!G@%�oMR ubj�  h)��}�(h G@N���v�h!G@48�ubj�  h)��}�(h G@N��>�bh!G@3ό�ݚ�ubj�  h)��}�(h G@@���eh!G@"�Ó��ubj�  hA)��}�(hDG��
 � � hEG��|��FhFG?�����ubj�  G@F�ZROj�  G?֦�)O]j�  G@=��'�ǧubj�  Kj�  �j�  hubj�  hj�  h)��}�(h G���,�<�`h!G��l��}Ӏubj�  h)��}�(h G��t?�լ h!G?�U�ٺ� ubj�  Kj�  �j�  h)��}�(h G        h!G        ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(h,j�  j�  hj�  h)��}�(h G?�*Z\mTh!G?�Oc.�hubj�  h)��}�(h G��t?�լ h!G?�U�ٺ� ubj�  Kj�  �j�  h)��}�(h G@-Kك�_�h!G@ ��z��ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(h,j�  j�  hj�  h)��}�(h G@;�R#Nh!G@%�oMR ubj�  h)��}�(h G��t?�լ h!G?�U�ٺ� ubj�  Kj�  �j�  h)��}�(h G@, ���z\h!G@y�8K/�ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(h,j�  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G@>A\L��Nh!G@0���ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG@F�ZROubj�  j�  )��}�(j�  h)��}�(h K h!K ubj�  h)��}�(h G@O5�ԍ|h!G@C���̖�ubj�  h)��}�(h G@]��x�h!G@L�Xp-ubj�  h)��}�(h G@]��x�h!G@L�Xp-ubj�  h)��}�(h G@Ln	Xc4h!G@2$����ubj�  hA)��}�(hDG��(�!ѵxhEG��_��fhFG?���|,�!ubj�  G?�������j�  G?�g���j�  G@Rv��u�ubj�  Kj�  �j�  hubj�  hj�  h)��}�(h G@O5�ԍ|h!G@C���̖�ubj�  h)��}�(h K h!K ubj�  Kj�  �j�  h)��}�(h G@>A\L��Nh!G@0���ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G@F�ZROubjZ  )��}�(j5  j8  )��}�(j;  hj<  j�  j=  Nj>  j�  j?  K hh)��}�(hhj�  j�  j�  j�  j�  j�  ububhjC  j]  j�  j^  jH  j�  hubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j  ubjZ  )��}�(j5  jA  hjC  j]  j/  j^  j�  j�  hubj`  )��}�(j]  j/  jc  jK  ubj`  )��}�(j]  j/  jc  jQ  ubj`  )��}�(j]  j/  jc  jW  ubj`  )��}�(j]  j/  jc  j]  ubj`  )��}�(j]  j/  jc  jc  ubj`  )��}�(j]  j/  jc  ji  ubj`  )��}�(j]  j/  jc  jo  ubjZ  )��}�(j5  jA  hjC  j]  j�  j^  j/  j�  hubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubjZ  )��}�(j5  jA  hjC  j]  j  j^  j�  j�  hubj`  )��}�(j]  j  jc  j+  ubj`  )��}�(j]  j  jc  j1  ubj`  )��}�(j]  j  jc  j7  ubj`  )��}�(j]  j  jc  j=  ubjZ  )��}�(j5  jA  hjC  j]  jU  j^  j  j�  hubj`  )��}�(j]  jU  jc  jq  ubj`  )��}�(j]  jU  jc  jw  ubj`  )��}�(j]  jU  jc  j}  ubj`  )��}�(j]  jU  jc  j�  ubj`  )��}�(j]  jU  jc  j�  ubj`  )��}�(j]  jU  jc  j�  ubj`  )��}�(j]  jU  jc  j�  ubj`  )��}�(j]  jU  jc  j�  ubjZ  )��}�(j5  jA  hjC  j]  j�  j^  jU  j�  hubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubjZ  )��}�(j5  jA  hjC  j]  j�  j^  j�  j�  hubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j!  ubj`  )��}�(j]  j�  jc  j'  ubjZ  )��}�(j5  jA  hjC  j]  j?  j^  j�  j�  hubj`  )��}�(j]  j?  jc  j[  ubj`  )��}�(j]  j?  jc  ja  ubj`  )��}�(j]  j?  jc  jg  ubj`  )��}�(j]  j?  jc  jm  ubj`  )��}�(j]  j?  jc  js  ubj`  )��}�(j]  j?  jc  jy  ubj`  )��}�(j]  j?  jc  j  ubj`  )��}�(j]  j?  jc  j�  ubj`  )��}�(j]  j?  jc  j�  ubj`  )��}�(j]  j?  jc  j�  ubj`  )��}�(j]  j?  jc  j�  ubj`  )��}�(j]  j?  jc  j�  ubjZ  )��}�(j5  jA  hjC  j]  j�  j^  j?  j�  hubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubjZ  )��}�(j5  jA  hjC  j]  j  j^  j�  j�  hubj`  )��}�(j]  j  jc  j/  ubj`  )��}�(j]  j  jc  j5  ubj`  )��}�(j]  j  jc  j;  ubj`  )��}�(j]  j  jc  jA  ubjZ  )��}�(j5  jA  hjC  j]  jY  j^  j  j�  hubj`  )��}�(j]  jY  jc  ju  ubj`  )��}�(j]  jY  jc  j{  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubj`  )��}�(j]  jY  jc  j�  ubjZ  )��}�(j5  jA  hjC  j]  j�  j^  jY  j�  hubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j	  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j  ubj`  )��}�(j]  j�  jc  j!  ubj`  )��}�(j]  j�  jc  j'  ubj`  )��}�(j]  j�  jc  j-  ubj`  )��}�(j]  j�  jc  j3  ubj`  )��}�(j]  j�  jc  j9  ubj`  )��}�(j]  j�  jc  j?  ubj`  )��}�(j]  j�  jc  jE  ubj`  )��}�(j]  j�  jc  jK  ubj`  )��}�(j]  j�  jc  jQ  ubj`  )��}�(j]  j�  jc  jW  ubj`  )��}�(j]  j�  jc  j]  ubj`  )��}�(j]  j�  jc  jc  ubj`  )��}�(j]  j�  jc  ji  ubj`  )��}�(j]  j�  jc  jo  ubj`  )��}�(j]  j�  jc  ju  ubj`  )��}�(j]  j�  jc  j{  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj`  )��}�(j]  j�  jc  j�  ubj�  )��}�(h,j�  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G@K"/�i"�h!G@>�-��ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG@������ubj�  j�  )��}�(j�  h)��}�(h K h!K ubj�  h)��}�(h G@S��̝�Nh!G@;��M��jubj�  h)��}�(h G@`�f�?C
h!G@H<("��ubj�  h)��}�(h G@`�f�?C
h!G@H<("��ubj�  h)��}�(h G@K�����h!G@4Z�P��ubj�  hA)��}�(hDG?yĤ�H� hEG?yę����hFG?��ր$ubj�  G?�D�ôX%j�  G?գ^HxBj�  G@T�
��ubj�  Kj�  �j�  hubj�  hj�  h)��}�(h G@S��̝�Nh!G@;��M��jubj�  h)��}�(h K h!K ubj�  Kj�  �j�  h)��}�(h G@K"/�i"�h!G@>�-��ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G@������ube�version��0.0.1�u.