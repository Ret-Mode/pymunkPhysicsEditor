��~b      }�(�database��editorCode.database��Database���)��}�(�bodies�]�(�$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��BODY��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G?�N��>�h!G?��oPubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�51{  h!G?�Aw��|ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]�(�%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�N��>�h!G?�����ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�51{  h!G?�wJ_��ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��
elasticity�G        �friction�G?�      �isSensor���shapeFilterGroup�K �shapeFilterCategory������ �shapeFilterMask������ �type��Polygon��internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G@Ҙ���h!G���x4���ubh"h)��}�(h G@Ҙ���h!G���x4���ububh)��}�(hh)��}�(h G?䪘���h!G��#��u�ubh"h)��}�(h G?䪘���h!G��#��u�ububh)��}�(hh)��}�(h G�����0h!G���7�E�ubh"h)��}�(h G�����0h!G���7�E�ububh)��}�(hh)��}�(h G����h�Uh!G?�*��R� ubh"h)��}�(h G����h�Uh!G?�*��R� ububh)��}�(hh)��}�(h G�	��]"�h!G?���ah�(ubh"h)��}�(h G�	��]"�h!G?���ah�(ububh)��}�(hh)��}�(h G@�u9��h!G?�����{\ubh"h)��}�(h G@�u9��h!G?�����{\ububh)��}�(hh)��}�(h G@������h!G?ǟ�}]0�ubh"h)��}�(h G@������h!G?ǟ�}]0�ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G�H��sUsh!G?�"֩$sub�user�h)��}�(h G        h!G        ubh"h)��}�(h G�H��sUsh!G?�"֩$sub�userDefined��ub�area�G@�ˠ�%��density�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h��ub�mass�h�)��}�(h�G?�      h�G        h"G@�ˠ�%�h��ub�moment�h�)��}�(h�G@4I��#�#h�G        h"G@4I��#�#h��ubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G��s��-�h!G?�U�����ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�,!��Lh!G?ϳ�"��ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1�hfG        hgG?�      hh�hiK hj����� hk����� hlhmhnhq)��}�(ht]�(h)��}�(hh)��}�(h G���Gp�h!G?����Subh"h)��}�(h G���Gp�h!G?����Sububh)��}�(hh)��}�(h G���#���h!G?�P�LUubh"h)��}�(h G���#���h!G?�P�LUububh)��}�(hh)��}�(h G?��ՠ�� h!G?���ubh"h)��}�(h G?��ՠ�� h!G?���ububh)��}�(hh)��}�(h G?��_j"-�h!G?�h��C0ubh"h)��}�(h G?��_j"-�h!G?�h��C0ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G��st���h!G?��Z����ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��st���h!G?��Z����ubh��ubh�G?��/r�b�h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G?��/r�b�h��ubh�h�)��}�(h�G?�=(lh�G        h"G?�=(lh��ubububehl�Dynamic�h��+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G��</"*�h!G?�{A�0ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��</"*�h!G?�{A�0ubh��ubh�G@=}�~@h�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@=}�~@h�G@r�     h"G@r�     h��ubh�h�)��}�(h�G@5�����dh�G        h"G@5�����dh��ubububh)��}�(h�Wheel�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G������?0h!G��g���ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G������?0h9G        h:G?�      h;G��g���ubh<h)��}�(h G������?0h!G��g���ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�hJ�Circle���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G������?0h!G��g���ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G������?0h9G        h:G?�      h;G��g���ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfG        hgG@4      hh�hiK hj����� hk����� hl�Circle�hnho�
CircleSpec���)��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj[  �radiusVector�h)��}�(h G        h!G        ubh�h�CircleRadius���)��}�(h"G?�      �base�G?�      ub�	drawLines�K ubh�h��CirclePhysics���)��}�(h�h�)��}�(h�h)��}�(h G������?0h!G��g���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububahlj  h�j  )��}�(h�h�)��}�(h�h)��}�(h G������?0h!G��g���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@	!�TD-h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububh)��}�(h�Wheel2�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G@ϔ��ph9G        h:G?�      h;G��Ù���<ubh<h)��}�(h G@ϔ��ph!G��Ù���<ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�j;  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G@ϔ��ph9G        h:G?�      h;G��Ù���<ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hfG        hgG@4      hh�hiK hj����� hk����� hljU  hnjW  )��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj�  jg  h)��}�(h G        h!G        ubh�jk  )��}�(h"G?�      jn  G?�      ubjo  K ubh�jq  )��}�(h�h�)��}�(h�h)��}�(h G@ϔ��ph!G��Ù���<ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububahlj  h�j  )��}�(h�h�)��}�(h�h)��}�(h G@ϔ��ph!G��Ù���<ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@	!�TD-h�G@r�     h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ububube�	shapeList�]�(hMh�j<  j�  e�constraints�]�(�/editorCode.constraintInternals.editorConstraint��GrooveJoint���)��}�(h�CNSTRNT�hl�Groove��bodyA�h�bodyB�j   �selfCollide���maxForce�G�      �maxBias�G�      �	errorBias�G?]q5�NZ�grooveA�h�OffsetPoint���)��}�(�offset�h)��}�(h G��u�Şbh!G��F�!$��ubhh)��}�(h G��u�Şbh!G��F�!$��ubh"h)��}�(h G������?0h!G��g���ubub�grooveB�j  )��}�(j  h)��}�(h G��GGw@"h!G?��x��r ubhh)��}�(h G��GGw@"h!G?��x��r ubh"h)��}�(h G���	����h!G?�\X�I0ubub�anchorB�j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububj�  )��}�(h�	CNSTRNT_1�hlj  j  hj  j�  j  �j  G�      j  G�      j  G?]q5�NZj	  j  )��}�(j  h)��}�(h G@ݱ��h!G���`�*Hubhh)��}�(h G@ݱ��h!G���`�*Hubh"h)��}�(h G@ϔ��ph!G��Ù���<ububj  j  )��}�(j  h)��}�(h G@ݱ��h!G���qv� ubhh)��}�(h G@ݱ��h!G���qv� ubh"h)��}�(h G@ϔ��ph!G?�����ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubububj�  �DampedSpring���)��}�(h�	CNSTRNT_2�hl�Damped Spring�j  hj  j   j  �j  G�      j  G�      j  G?]q5�NZ�
restLength�G        �	stiffness�G@@     �damping�G?�      �anchorA�j  )��}�(j  h)��}�(h G��u�Şbh!G��F�!$��ubhh)��}�(h G��u�Şbh!G��F�!$��ubh"h)��}�(h G������?0h!G��g���ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububjC  )��}�(h�	CNSTRNT_3�hljG  j  hj  j�  j  �j  G�      j  G�      j  G?]q5�NZjH  G        jI  G@@     jJ  G?�      jK  j  )��}�(j  h)��}�(h G@ݱ��h!G���`�*Hubhh)��}�(h G@ݱ��h!G���`�*Hubh"h)��}�(h G@ϔ��ph!G��Ù���<ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububube�mappings�]�(�editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�      h!G��      ubh"h)��}�(h G�      h!G��      ububh)��}�(hh)��}�(h G@      h!G��      ubh"h)��}�(h G@      h!G��      ububh)��}�(hh)��}�(h G�      h!G?�      ubh"h)��}�(h G�      h!G?�      ububh)��}�(hh)��}�(h G@      h!G?�      ubh"h)��}�(h G@      h!G?�      ubube�textureSize�]�(M K`e�anchor�]�(G@`      G@H      e�mappingSize�]�(M K`e�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@`      h!G@H      ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububjs  )��}�(h�MAP:1�jw  Kjx  j   h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G������?0h9G        h:G?�      h;G��g���ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G�|��t�h!G�3��Y�tububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G���OI�~`h!G�3��Y�tububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G�|��t�h!G�џ�B��ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G���OI�~`h!G�џ�B��ububej�  ]�(K@K@ej�  ]�(G@@      G@@      ej�  ]�(K@K@ej�  ]�(K K ej�  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububjs  )��}�(h�MAP:1_1�jw  Kjx  j�  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G@ϔ��ph9G        h:G?�      h;G��Ù���<ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?�7�)��h!G� a��I�ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@
ϔ��ph!G� a��I�ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G?�7�)��h!G��s0�tǀububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G@
ϔ��ph!G��s0�tǀububej�  ]�(K@K@ej�  ]�(G@@      G@@      ej�  ]�(K@K@ej�  ]�(K K ej�  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubububeub�textureSizes�]�(M K`��K@K@��K K ��j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  e�texturePaths�]�(�data/textures/shark.png��data/textures/wheel1.png�� �j1  j1  j1  j1  j1  j1  j1  j1  j1  j1  j1  j1  j1  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�j�  �currentShape�j�  �currentConstraint�j\  �currentMapping�j�  �currentMappingChannel�Khh)��}�(hhj�  j�  j�  j�  jo  jp  ub�pivot�h)��}�(h G@ϔ��ph!G?�����ububhjH  �object�h�prevCurrent�Nubj:  )��}�(j=  jA  hjH  jM  j   jN  hubj:  )��}�(j=  jA  hjH  jM  j�  jN  j   ubj8  �ComSetBodyAsCurrent���)��}�(j=  jA  h�BODY_1��prev�j�  ubj8  �ComResetUserParam���)��}�(�param�j�  �oldUserFlag��ubjZ  )��}�(j]  j�  j^  �ubjZ  )��}�(j]  j�  j^  �ubj8  �ComResetUserCoords���)��}�(�coords�j�  j^  �ubj8  �ComRenameBody���)��}�(jx  j   hjH  �newName�j"  �oldName�jW  ubjT  )��}�(j=  jA  h�BODY_2�jX  j   ubjZ  )��}�(j]  j�  j^  �ubjZ  )��}�(j]  j�  j^  �ubjZ  )��}�(j]  j�  j^  �ubjd  )��}�(jg  j�  j^  �ubji  )��}�(jx  j�  hjH  jl  j�  jm  jp  ubjT  )��}�(j=  jA  hhjX  j�  ubj8  �ComLoadTexture���)��}�(hjH  �newPath�j/  �destChannel�K �newSize�j*  �oldPath�j1  �oldSize�j,  ubj~  )��}�(hjH  j�  j0  j�  Kj�  K@K@��j�  j1  j�  j,  ubj~  )��}�(hjH  j�  j0  j�  Kj�  j+  j�  j0  j�  j�  ubj8  �ComCreateMapping���)��}�(j=  jA  hjH  �mapping�jt  �prevMapping�Nubj�  )��}�(j=  jA  hjH  j�  j�  j�  Nubj�  )��}�(j=  jA  hjH  j�  j�  j�  j�  ubj8  �ComAddNewShape���)��}�(j=  jA  hjH  �shape�hM�	prevShape�Njx  hubj8  �ComNewShapeAddPoint���)��}�(j�  hM�point�hvubj�  )��}�(j�  hMj�  h|ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j=  jA  hjH  j�  h�j�  hMjx  hubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj8  �ComSelectNextBody���)��}�(j=  jA  �oldBody�h�oldShape�hƌnewBody�j   �newShape�N�executed��ubj8  �ComSelectPrevBody���)��}�(j=  jA  j�  j   j�  j;  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G        h!G        ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfG        hgG?�      hh�hiK hj����� hk����� hljU  hnjW  )��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj�  jg  h)��}�(h G        h!G        ubh�jk  )��}�(h"G?�      jn  G?�      ubjo  K ubh�jq  )��}�(h�h�)��}�(h�h)��}�(h G        h!G        ubh�h)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububj�  hj�  h�j�  �ubj�  )��}�(j=  jA  j�  hj�  h�j�  j   j�  Nj�  �ubj�  )��}�(j=  jA  hjH  j�  j<  j�  Njx  j   ubj�  )��}�(j=  jA  j�  j   j�  j<  j�  j�  j�  Nj�  �ubj�  )��}�(j=  jA  hjH  j�  j�  j�  Njx  j�  ubj�  )��}�(j=  jA  j�  j�  j�  j�  j�  j   j�  j<  j�  �ubj�  )��}�(j=  jA  j�  j   j�  j<  j�  j�  j�  j�  j�  �ubj8  �ComSetMappingFromSelection���)��}�(j�  j�  �	selection�h�	Selection���)��}�(�start�h)��}�(h G@_@i��h!G�A"\���ub�end�h)��}�(h G�@w9e��h!G@V�&7kM0ub�active��ub�	oldOffset�j  j�  j  ubj  )��}�(j�  j�  j  j  j  j  j�  j  ubj8  �ComSetPivot���)��}�(jJ  jK  �newWorld�h)��}�(h G������?0h!G��g���ub�oldWorld�h)��}�(h G        h!G        ububjT  )��}�(j=  jA  hj"  jX  j�  ubj8  �ComMoveObject���)��}�(�obj�j   �forward�h)��}�(h G������?0h!G��g���ububj  )��}�(jJ  jK  j"  h)��}�(h G@ϔ��ph!G��Ù���<ubj%  h)��}�(h G������?0h!G��g���ububjT  )��}�(j=  jA  hj�  jX  j   ubj+  )��}�(j.  j�  j/  h)��}�(h G@ϔ��ph!G��Ù���<ububj8  �ComAddConstraint���)��}�(hjH  j=  jA  jM  j�  jN  Nubj8  �ComConstraintSetNewBodyA���)��}�(�entity�j�  j�  hj�  Nubj8  �ComConstraintSetNewBodyB���)��}�(jF  j�  j�  j   j�  Nubj8  �ComSetGrooveAFromCoords���)��}�(jF  j�  �	newXValue�G��u�Şb�	newYValue�G��F�!$��	oldXValue�G        �	oldYValue�G        ubj  )��}�(jJ  jK  j"  h)��}�(h G���	����h!G?�\X�I0ubj%  h)��}�(h G@ϔ��ph!G��Ù���<ububj8  �ComSetGrooveBFromCoords���)��}�(jF  j�  jO  G��GGw@"jP  G?��x��r jQ  G        jR  G        ubj?  )��}�(hjH  j=  jA  jM  j'  jN  j�  ubj8  �ComSetConstraintAsCurrent���)��}�(j=  jA  hj)  jX  j'  ubjC  )��}�(jF  j'  j�  hj�  NubjH  )��}�(jF  j'  j�  j   j�  NubjH  )��}�(jF  j'  j�  j�  j�  j   ubjL  )��}�(jF  j'  jO  G@ݱ��jP  G���`�*HjQ  G        jR  G        ubj  )��}�(jJ  jK  j"  h)��}�(h G@ϔ��ph!G?�����ubj%  h)��}�(h G���	����h!G?�\X�I0ububjZ  )��}�(jF  j'  jO  G@ݱ��jP  G���qv� jQ  G        jR  G        ubj?  )��}�(hjH  j=  jA  jM  jD  jN  j'  ubjC  )��}�(jF  jD  j�  hj�  NubjH  )��}�(jF  jD  j�  j   j�  Nubj8  �ComSetAnchorAFromCoords���)��}�(jF  jD  jO  G        jP  G        jQ  G        jR  G        ubjz  )��}�(jF  jD  jO  G��u�ŞbjP  G��F�!$��jQ  G        jR  G        ubj8  �ComSetRestLength���)��}�(jF  jD  �newValue�G        �oldValue�G?�      ubj`  )��}�(j=  jA  hjF  jX  jD  ubj8  �ComConstraintClone���)��}�(hjH  j=  jA  �baseConstraint�jD  �newConstraint�j\  �index�Kubj`  )��}�(j=  jA  hj^  jX  j\  ubjH  )��}�(jF  j\  j�  j�  j�  j   ubjz  )��}�(jF  j\  jO  G@ݱ��jP  G���`�*HjQ  G��u�ŞbjR  G��F�!$��ubjT  )��}�(j=  j@  )��}�(jC  hjD  h�jE  j\  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhhjX  j�  ubjT  )��}�(j=  j�  hj"  jX  hubjT  )��}�(j=  j�  hj�  jX  j   ubjT  )��}�(j=  j�  hhjX  j�  ubj`  )��}�(j=  j�  hjF  jX  j\  ubj8  �ComSetStiffness���)��}�(jF  jD  j�  G@�@     j�  G?�      ubj8  �ComSetDamping���)��}�(jF  jD  j�  G@I      j�  G?�      ubj`  )��}�(j=  j�  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@�@     j�  G?�      ubj�  )��}�(jF  j\  j�  G@I      j�  G?�      ubj`  )��}�(j=  j@  )��}�(jC  j�  jD  j�  jE  jD  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhjF  jX  j\  ubj8  �ComSetUserParam���)��}�(j]  j�  j^  ��
oldUserVal�G        �value�G@r�     ubjT  )��}�(j=  j@  )��}�(jC  j�  jD  j�  jE  j\  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhhjX  j�  ubj�  )��}�(j=  j�  j�  hj�  h�j�  j   j�  j<  j�  �ubj8  �ComNewShapeSetFriction���)��}�(j�  j<  j�  G?�      j�  G@4      ubj�  )��}�(j=  j�  j�  j   j�  j<  j�  j�  j�  j�  j�  �ubj�  )��}�(j�  j�  j�  G?�      j�  G@4      ubj`  )��}�(j=  j@  )��}�(jC  j�  jD  j�  jE  j\  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@i      j�  G@�@     ubj�  )��}�(jF  jD  j�  G@Y      j�  G@I      ubj`  )��}�(j=  j�  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@i      j�  G@�@     ubj�  )��}�(jF  j\  j�  G@Y      j�  G@I      ubj`  )��}�(j=  j@  )��}�(jC  j�  jD  j�  jE  j\  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jF  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jF  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jF  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jF  jD  j�  G@È     j�  G@i      ubj�  )��}�(jF  jD  j�  G@Y      j�  G@Y      ubj`  )��}�(j=  j�  hj^  jX  jD  ubj`  )��}�(j=  j�  hjF  jX  j\  ubj`  )��}�(j=  j�  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@È     j�  G@i      ubj�  )��}�(jF  j\  j�  G@Y      j�  G@Y      ubj�  )��}�(jF  j\  j�  G@Y      j�  G@Y      ubj�  )��}�(jF  j\  j�  G@Y      j�  G@Y      ubj`  )��}�(j=  j@  )��}�(jC  j�  jD  j�  jE  j\  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@�@     j�  G@È     ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@�@     j�  G@È     ubj`  )��}�(j=  j@  )��}�(jC  j�  jD  j�  jE  j\  jF  j�  jG  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubjJ  h)��}�(h G        h!G        ububhjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@I      j�  G@Y      ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@I      j�  G@Y      ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(hj  j=  j  j�  jD  j�  jC  )��}�(h�	CNSTRNT_4�hl�Damped Spring�j  hj  j   j  �j  G�      j  G�      j  G?]q5�NZjH  G        jI  G@�@     jJ  G@I      jK  j  )��}�(j  h)��}�(h G��u�Şbh!G��F�!$��ubhh)��}�(h G��u�Şbh!G��F�!$��ubh"h)��}�(h G������?0h!G��g���ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububj�  Kubj`  )��}�(j=  j  hj(  jX  j&  ubj`  )��}�(j=  j  hjF  jX  j&  ubj`  )��}�(j=  j  hj(  jX  jD  ubj`  )��}�(j=  j  hj^  jX  j&  ubj�  )��}�(hj  j=  j  j�  j\  j�  jC  )��}�(h�	CNSTRNT_5�hlj)  j  hj  j�  j  �j  G�      j  G�      j  G?]q5�NZjH  G        jI  G@�@     jJ  G@I      jK  j  )��}�(j  h)��}�(h G@ݱ��h!G���`�*Hubhh)��}�(h G@ݱ��h!G���`�*Hubh"h)��}�(h G@ϔ��ph!G��Ù���<ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubububj�  Kubj`  )��}�(j=  j  hjF  jX  jD  ubj8  �ComDelConstraint���)��}�(hj  j=  j  jM  jD  �objIndex�Kubj`  )��}�(j=  j  hj(  jX  j\  ubjZ  )��}�(hj  j=  j  jM  j&  j]  Kubj�  )��}�(jF  j\  j�  G@�@     j�  G@I      ubj�  )��}�(jF  j\  j�  G@Y      j�  G@�@     ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@Y      j�  G@�@     ubj�  )��}�(jF  jD  j�  G@�@     j�  G@I      ubj�  )��}�(jF  jD  j�  G@$      j�  G@Y      ubj�  )��}�(jF  jD  j�  G@È     j�  G@�@     ubj`  )��}�(j=  j  hj^  jX  jD  ubj`  )��}�(j=  j  hjF  jX  j\  ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@$      j�  G@Y      ubj�  )��}�(jF  j\  j�  G@È     j�  G@�@     ubj�  )��}�(jF  j\  j�  G@@     j�  G@$      ubj`  )��}�(j=  j  hj^  jX  j\  ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@@     j�  G@$      ubj�  )��}�(jF  jD  j�  G@@     j�  G@È     ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@@     j�  G@È     ubj`  )��}�(j=  j  hj^  jX  j\  ubj`  )��}�(j=  j  hjF  jX  j\  ubj`  )��}�(j=  j  hj^  jX  jD  ubj`  )��}�(j=  j  hjF  jX  j\  ubj`  )��}�(j=  j  hj^  jX  jD  ubj`  )��}�(j=  j  hjF  jX  j\  ubj`  )��}�(j=  j  hjF  jX  jD  ubj�  )��}�(jF  jD  j�  G@4      j�  G@@     ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@4      j�  G@@     ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@4      j�  G@@     ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@4      j�  G@@     ubj�  )��}�(jF  j\  j�  G@i      j�  G@4      ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@i      j�  G@4      ubj`  )��}�(j=  j  hjF  jX  jD  ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G?�      j�  G@4      ubj`  )��}�(j=  j  hj^  jX  j\  ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G?�      j�  G@4      ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@È     j�  G@i      ubj`  )��}�(j=  j  hj^  jX  j\  ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@È     j�  G@i      ubj�  )��}�(jF  jD  j�  G@��     j�  G@È     ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@��     j�  G@È     ubj�  )��}�(jF  j\  j�  G@��     j�  G@��     ubj`  )��}�(j=  j  hjF  jX  j\  ubj�  )��}�(jF  jD  j�  G@��     j�  G@��     ubj�  )��}�(jF  jD  j�  G@@     j�  G@��     ubj`  )��}�(j=  j  hjF  jX  jD  ubj`  )��}�(j=  j  hj^  jX  jD  ubj�  )��}�(jF  j\  j�  G@@     j�  G@��     ubjT  )��}�(j=  j@  )��}�(jC  hjD  h�jE  j\  jF  j�  jG  KhhjJ  h)��}�(h G        h!G        ububhj�  jX  j�  ubjZ  )��}�(j]  j�  j^  �ubjT  )��}�(j=  j�  hj"  jX  j�  ubjT  )��}�(j=  j�  hhjX  j   ubj�  )��}�(j]  j  j^  �j�  G        j�  G@r�     ube�version��0.0.2�u.