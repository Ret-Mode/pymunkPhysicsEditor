��4m      }�(�database��editorCode.database��Database���)��}�(�bodies�]�(�$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��BODY��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G?�N��>�h!G?��oPubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�51{  h!G?�Aw��|ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]�(�%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�N��>�h!G?�����ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�51{  h!G?�wJ_��ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��
elasticity�G        �friction�G?�      �isSensor���shapeFilterGroup�K �shapeFilterCategory������ �shapeFilterMask������ �type��Polygon��internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G@Ҙ���h!G���x4���ubh"h)��}�(h G@Ҙ���h!G���x4���ububh)��}�(hh)��}�(h G?䪘���h!G��#��u�ubh"h)��}�(h G?䪘���h!G��#��u�ububh)��}�(hh)��}�(h G�����0h!G���7�E�ubh"h)��}�(h G�����0h!G���7�E�ububh)��}�(hh)��}�(h G����h�Uh!G?�*��R� ubh"h)��}�(h G����h�Uh!G?�*��R� ububh)��}�(hh)��}�(h G�	��]"�h!G?���ah�(ubh"h)��}�(h G�	��]"�h!G?���ah�(ububh)��}�(hh)��}�(h G@�u9��h!G?�����{\ubh"h)��}�(h G@�u9��h!G?�����{\ububh)��}�(hh)��}�(h G@������h!G?ǟ�}]0�ubh"h)��}�(h G@������h!G?ǟ�}]0�ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G�H��sUsh!G?�"֩$sub�user�h)��}�(h G        h!G        ubh"h)��}�(h G�H��sUsh!G?�"֩$sub�userDefined��ub�area�G@�ˠ�%��density�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h��ub�mass�h�)��}�(h�G?�      h�G        h"G@�ˠ�%�h��ub�moment�h�)��}�(h�G@4I��#�#h�G        h"G@4I��#�#h��ubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G��s��-�h!G?�U�����ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�,!��Lh!G?ϳ�"��ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1�hfG        hgG?�      hh�hiK hj����� hk����� hlhmhnhq)��}�(ht]�(h)��}�(hh)��}�(h G���Gp�h!G?����Subh"h)��}�(h G���Gp�h!G?����Sububh)��}�(hh)��}�(h G���#���h!G?�P�LUubh"h)��}�(h G���#���h!G?�P�LUububh)��}�(hh)��}�(h G?��ՠ�� h!G?���ubh"h)��}�(h G?��ՠ�� h!G?���ububh)��}�(hh)��}�(h G?��_j"-�h!G?�h��C0ubh"h)��}�(h G?��_j"-�h!G?�h��C0ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G��st���h!G?��Z����ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��st���h!G?��Z����ubh��ubh�G?��/r�b�h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G?��/r�b�h��ubh�h�)��}�(h�G?�=(lh�G        h"G?�=(lh��ubububehl�Dynamic�h��+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G��</"*�h!G?�{A�0ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��</"*�h!G?�{A�0ubh��ubh�G@=}�~@h�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@=}�~@h�G@��     h"G@��     h��ubh�h�)��}�(h�G@5�����dh�G@i      h"G@i      h��ubububh)��}�(h�Wheel�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G������?0h!G��g���ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G������?0h9G        h:G?�      h;G��g���ubh<h)��}�(h G������?0h!G��g���ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�hJ�Circle���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G������?0h!G��g���ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G������?0h9G        h:G?�      h;G��g���ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfG        hgG@4      hh�hiK hj����� hk����� hl�Circle�hnho�
CircleSpec���)��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj[  �radiusVector�h)��}�(h G        h!G        ubh�h�CircleRadius���)��}�(h"G?�      �base�G?�      ub�	drawLines�K ubh�h��CirclePhysics���)��}�(h�h�)��}�(h�h)��}�(h G������?0h!G��g���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububahlj  h�j  )��}�(h�h�)��}�(h�h)��}�(h G������?0h!G��g���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@	!�TD-h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububh)��}�(h�Wheel2�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G@ϔ��ph9G        h:G?�      h;G��Ù���<ubh<h)��}�(h G@ϔ��ph!G��Ù���<ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�j;  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G@ϔ��ph9G        h:G?�      h;G��Ù���<ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hfG        hgG@4      hh�hiK hj����� hk����� hljU  hnjW  )��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj�  jg  h)��}�(h G        h!G        ubh�jk  )��}�(h"G?�      jn  G?�      ubjo  K ubh�jq  )��}�(h�h�)��}�(h�h)��}�(h G@ϔ��ph!G��Ù���<ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ubububahlj  h�j  )��}�(h�h�)��}�(h�h)��}�(h G@ϔ��ph!G��Ù���<ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@	!�TD-h�G@r�     h"G@	!�TD-h��ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h��ububube�	shapeList�]�(hMh�j<  j�  e�constraints�]�(�/editorCode.constraintInternals.editorConstraint��GrooveJoint���)��}�(h�CNSTRNT�hl�Groove��bodyA�h�bodyB�j   �selfCollide���maxForce�G�      �maxBias�G�      �	errorBias�G?]q5�NZ�grooveA�h�OffsetPoint���)��}�(�offset�h)��}�(h G��u�Şbh!G��F�!$��ubhh)��}�(h G��u�Şbh!G��F�!$��ubh"h)��}�(h G������?0h!G��g���ubub�grooveB�j  )��}�(j  h)��}�(h G��GGw@"h!G?��x��r ubhh)��}�(h G��GGw@"h!G?��x��r ubh"h)��}�(h G���	����h!G?�\X�I0ubub�anchorB�j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububj�  )��}�(h�	CNSTRNT_1�hlj  j  hj  j�  j  �j  G�      j  G�      j  G?]q5�NZj	  j  )��}�(j  h)��}�(h G@ݱ��h!G���`�*Hubhh)��}�(h G@ݱ��h!G���`�*Hubh"h)��}�(h G@ϔ��ph!G��Ù���<ububj  j  )��}�(j  h)��}�(h G@ݱ��h!G���qv� ubhh)��}�(h G@ݱ��h!G���qv� ubh"h)��}�(h G@ϔ��ph!G?�����ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubububj�  �DampedSpring���)��}�(h�	CNSTRNT_2�hl�Damped Spring�j  hj  j   j  �j  G�      j  G�      j  G?]q5�NZ�
restLength�G        �	stiffness�G@�@     �damping�G@o@     �anchorA�j  )��}�(j  h)��}�(h G��u�Şbh!G��F�!$��ubhh)��}�(h G��u�Şbh!G��F�!$��ubh"h)��}�(h G������?0h!G��g���ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububjC  )��}�(h�	CNSTRNT_3�hljG  j  hj  j�  j  �j  G�      j  G�      j  G?]q5�NZjH  G        jI  G@�@     jJ  G@o@     jK  j  )��}�(j  h)��}�(h G@ݱ��h!G���`�*Hubhh)��}�(h G@ݱ��h!G���`�*Hubh"h)��}�(h G@ϔ��ph!G��Ù���<ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ububube�mappings�]�(�editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�      h!G��      ubh"h)��}�(h G�      h!G��      ububh)��}�(hh)��}�(h G@      h!G��      ubh"h)��}�(h G@      h!G��      ububh)��}�(hh)��}�(h G�      h!G?�      ubh"h)��}�(h G�      h!G?�      ububh)��}�(hh)��}�(h G@      h!G?�      ubh"h)��}�(h G@      h!G?�      ubube�textureSize�]�(M K`e�anchor�]�(G@`      G@H      e�mappingSize�]�(M K`e�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@_>�h!G@L��q�ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububjs  )��}�(h�MAP:1�jw  Kjx  j   h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G������?0h9G        h:G?�      h;G��g���ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G�|��t�h!G�3��Y�tububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G���OI�~`h!G�3��Y�tububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G�|��t�h!G�џ�B��ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G���OI�~`h!G�џ�B��ububej�  ]�(K@K@ej�  ]�(G@@      G@@      ej�  ]�(K@K@ej�  ]�(K K ej�  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububjs  )��}�(h�MAP:1_1�jw  Kjx  j�  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G@ϔ��ph9G        h:G?�      h;G��Ù���<ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?�7�)��h!G� a��I�ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@
ϔ��ph!G� a��I�ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G?�7�)��h!G��s0�tǀububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G@
ϔ��ph!G��s0�tǀububej�  ]�(K@K@ej�  ]�(G@@      G@@      ej�  ]�(K@K@ej�  ]�(K K ej�  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubububjs  )��}�(h�MAP:0_1�jw  K jx  hh,h.)��}�(h1h3)��}�(h6G@#ΝVj[�h7G        h8G�*]�<�?;h9G        h:G@#ΝVj[�h;G?�U��Ghubh<h)��}�(h G?�Lo�g2�h!G����5Loubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?��mѤ\ubj�  ]�(h)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G��Û2g��h!G?�X���ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G?�ٟzm'8h!G?�X���ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G��Û2g��h!G@�=-{�Vububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G?�ٟzm'8h!G@�=-{�Vububej�  ]�(M K`ej�  ]�(G@`      G@H      ej�  ]�(KK	ej�  ]�(K�K3ej�  ]�(h)��}�(h G?��     h!G?�      ubh)��}�(h G?��     h!G?�      ubh)��}�(h G?��     h!G?�      ubh)��}�(h G?��     h!G?�      ubeh�h)��}�(h G@eIR��|h!G@HMZ��ubj�  h)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G�ǧ����h!G@g��*�ubububeub�textureSizes�]�(M K`��K@K@��K K ��je  je  je  je  je  je  je  je  je  je  je  je  je  e�texturePaths�]�(�data/textures/shark.png��data/textures/wheel1.png�� �jj  jj  jj  jj  jj  jj  jj  jj  jj  jj  jj  jj  jj  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��ComConstraintSetNewBodyB���)��}�(�entity�jD  �newBody�j   �oldBody�Nubjq  �ComSetAnchorAFromCoords���)��}�(jv  jD  �	newXValue�G        �	newYValue�G        �	oldXValue�G        �	oldYValue�G        ubjz  )��}�(jv  jD  j}  G��u�Şbj~  G��F�!$��j  G        j�  G        ubjq  �ComSetRestLength���)��}�(jv  jD  �newValue�G        �oldValue�G?�      ubjq  �ComSetConstraintAsCurrent���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�j�  �currentShape�j�  �currentConstraint�j\  �currentMapping�j�  �currentMappingChannel�Khh)��}�(hhj�  j�  j�  j�  jo  jp  ub�pivot�h)��}�(h G@ϔ��ph!G?�����ububhjF  �prev�jD  ubjq  �ComConstraintClone���)��}�(hj�  j�  j�  �baseConstraint�jD  �newConstraint�j\  �index�Kubj�  )��}�(j�  j�  hj^  j�  j\  ubjs  )��}�(jv  j\  jw  j�  jx  j   ubjz  )��}�(jv  j\  j}  G@ݱ��j~  G���`�*Hj  G��u�Şbj�  G��F�!$��ubjq  �ComSetBodyAsCurrent���)��}�(j�  j�  )��}�(j�  hj�  h�j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhhj�  j�  ubj�  )��}�(j�  j�  hj"  j�  hubj�  )��}�(j�  j�  hj�  j�  j   ubj�  )��}�(j�  j�  hhj�  j�  ubj�  )��}�(j�  j�  hjF  j�  j\  ubjq  �ComSetStiffness���)��}�(jv  jD  j�  G@�@     j�  G?�      ubjq  �ComSetDamping���)��}�(jv  jD  j�  G@I      j�  G?�      ubj�  )��}�(j�  j�  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@�@     j�  G?�      ubj�  )��}�(jv  j\  j�  G@I      j�  G?�      ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  jD  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubjq  �ComSetUserParam���)��}�(�param�j�  �oldUserFlag���
oldUserVal�G        �value�G@r�     ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhhj�  j�  ubjq  �ComSelectNextBody���)��}�(j�  j�  jx  h�oldShape�h�jw  j   �newShape�j<  �executed��ubjq  �ComNewShapeSetFriction���)��}�(�shape�j<  j�  G?�      j�  G@4      ubj�  )��}�(j�  j�  jx  j   j�  j<  jw  j�  j�  j�  j�  �ubj�  )��}�(j�  j�  j�  G?�      j�  G@4      ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@i      j�  G@�@     ubj�  )��}�(jv  jD  j�  G@Y      j�  G@I      ubj�  )��}�(j�  j�  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@i      j�  G@�@     ubj�  )��}�(jv  j\  j�  G@Y      j�  G@I      ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jv  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jv  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jv  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(jv  jD  j�  G@È     j�  G@i      ubj�  )��}�(jv  jD  j�  G@Y      j�  G@Y      ubj�  )��}�(j�  j  hj^  j�  jD  ubj�  )��}�(j�  j  hjF  j�  j\  ubj�  )��}�(j�  j  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@È     j�  G@i      ubj�  )��}�(jv  j\  j�  G@Y      j�  G@Y      ubj�  )��}�(jv  j\  j�  G@Y      j�  G@Y      ubj�  )��}�(jv  j\  j�  G@Y      j�  G@Y      ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@�@     j�  G@È     ubj�  )��}�(j�  j)  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@�@     j�  G@È     ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@I      j�  G@Y      ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@I      j�  G@Y      ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(hj9  j�  j7  j�  jD  j�  jC  )��}�(h�	CNSTRNT_4�hl�Damped Spring�j  hj  j   j  �j  G�      j  G�      j  G?]q5�NZjH  G        jI  G@�@     jJ  G@I      jK  j  )��}�(j  h)��}�(h G��u�Şbh!G��F�!$��ubhh)��}�(h G��u�Şbh!G��F�!$��ubh"h)��}�(h G������?0h!G��g���ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G������?0h!G��g���ubububj�  Kubj�  )��}�(j�  j7  hjI  j�  jG  ubj�  )��}�(j�  j7  hjF  j�  jG  ubj�  )��}�(j�  j7  hjI  j�  jD  ubj�  )��}�(j�  j7  hj^  j�  jG  ubj�  )��}�(hj9  j�  j7  j�  j\  j�  jC  )��}�(h�	CNSTRNT_5�hljJ  j  hj  j�  j  �j  G�      j  G�      j  G?]q5�NZjH  G        jI  G@�@     jJ  G@I      jK  j  )��}�(j  h)��}�(h G@ݱ��h!G���`�*Hubhh)��}�(h G@ݱ��h!G���`�*Hubh"h)��}�(h G@ϔ��ph!G��Ù���<ububj  j  )��}�(j  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@ϔ��ph!G��Ù���<ubububj�  Kubj�  )��}�(j�  j7  hjg  j�  je  ubjq  �ComDelConstraint���)��}�(hj9  j�  j7  �object�je  �objIndex�Kubj�  )��}�(j�  j7  hjI  j�  j\  ubj{  )��}�(hj9  j�  j7  j~  jG  j  Kubj�  )��}�(jv  j\  j�  G@�@     j�  G@I      ubj�  )��}�(jv  j\  j�  G@Y      j�  G@�@     ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@Y      j�  G@�@     ubj�  )��}�(jv  jD  j�  G@�@     j�  G@I      ubj�  )��}�(jv  jD  j�  G@$      j�  G@Y      ubj�  )��}�(jv  jD  j�  G@È     j�  G@�@     ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@$      j�  G@Y      ubj�  )��}�(jv  j\  j�  G@È     j�  G@�@     ubj�  )��}�(jv  j\  j�  G@@     j�  G@$      ubj�  )��}�(j�  j7  hj^  j�  j\  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@@     j�  G@$      ubj�  )��}�(jv  jD  j�  G@@     j�  G@È     ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@@     j�  G@È     ubj�  )��}�(j�  j7  hj^  j�  j\  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(j�  j7  hjF  j�  jD  ubj�  )��}�(jv  jD  j�  G@4      j�  G@@     ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@4      j�  G@@     ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@4      j�  G@@     ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@4      j�  G@@     ubj�  )��}�(jv  j\  j�  G@i      j�  G@4      ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@i      j�  G@4      ubj�  )��}�(j�  j7  hjF  j�  jD  ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G?�      j�  G@4      ubj�  )��}�(j�  j7  hj^  j�  j\  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G?�      j�  G@4      ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@È     j�  G@i      ubj�  )��}�(j�  j7  hj^  j�  j\  ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@È     j�  G@i      ubj�  )��}�(jv  jD  j�  G@��     j�  G@È     ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@��     j�  G@È     ubj�  )��}�(jv  j\  j�  G@��     j�  G@��     ubj�  )��}�(j�  j7  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@��     j�  G@��     ubj�  )��}�(jv  jD  j�  G@@     j�  G@��     ubj�  )��}�(j�  j7  hjF  j�  jD  ubj�  )��}�(j�  j7  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@@     j�  G@��     ubj�  )��}�(j�  j�  )��}�(j�  hj�  h�j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhj�  j�  j�  ubjq  �ComResetUserParam���)��}�(j�  j�  j�  �ubj�  )��}�(j�  j�  hj"  j�  j�  ubj�  )��}�(j�  j�  hhj�  j   ubj�  )��}�(j�  j  j�  �j�  G        j�  G@r�     ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  j\  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@I      j�  G?�      ubj�  )��}�(j�  j
  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@I      j�  G?�      ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  jD  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhj^  j�  j\  ubj�  )��}�(jv  j\  j�  G@�@     j�  G@@     ubj�  )��}�(j�  j  hj^  j�  j\  ubj�  )��}�(j�  j  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@�@     j�  G@@     ubj�  )��}�(jv  j\  j�  G@@     j�  G@I      ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  jD  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@@     j�  G@I      ubj�  )��}�(j�  j*  hj^  j�  jD  ubj�  )��}�(j�  j*  hjF  j�  j\  ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  jD  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhj^  j�  j\  ubj�  )��}�(jv  j\  j�  G@I      j�  G@@     ubj�  )��}�(jv  j\  j�  G@�@     j�  G@�@     ubj�  )��}�(j�  j8  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@�@     j�  G@�@     ubj�  )��}�(jv  jD  j�  G@I      j�  G@@     ubj�  )��}�(j�  j�  )��}�(j�  j�  j�  j�  j�  jD  j�  j�  j�  Khh)��}�(hhj�  j�  j�  j�  jo  jp  ubj�  h)��}�(h G        h!G        ububhjF  j�  j\  ubj�  )��}�(j�  jJ  hj^  j�  jD  ubj�  )��}�(j�  jJ  hjF  j�  j\  ubj�  )��}�(j�  jJ  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@��     j�  G@�@     ubj�  )��}�(j�  jJ  hj^  j�  j\  ubj�  )��}�(j�  jJ  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@��     j�  G@�@     ubj�  )��}�(j�  j�  )��}�(j�  hj�  h�j�  j\  j�  j(  j�  K hhj�  h)��}�(h G?�ۂ�Wz�h!G?՜�5�E�ububhjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@Y      j�  G@I      ubj�  )��}�(j�  j`  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@Y      j�  G@I      ubj�  )��}�(j�  j`  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@b�     j�  G@Y      ubj�  )��}�(j�  j`  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@b�     j�  G@Y      ubj�  )��}�(j�  j`  hhj�  j�  ubj�  )��}�(j�  j  j�  �j�  G@r�     j�  G@��     ubj�  )��}�(jv  j\  j�  G@�X     j�  G@��     ubj�  )��}�(j�  j`  hj^  j�  j\  ubj�  )��}�(j�  j`  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@�X     j�  G@��     ubj�  )��}�(jv  jD  j�  G@i      j�  G@b�     ubj�  )��}�(j�  j`  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@i      j�  G@b�     ubj�  )��}�(j�  j`  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@�@     j�  G@�X     ubj�  )��}�(j�  j`  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@�@     j�  G@�X     ubj�  )��}�(j�  j`  hhj�  hubj�  )��}�(j�  j`  hj"  j�  hubjq  �ComStartTransform���)��}�(h,�editorCode.editorViewTransform��ContinuousTransform���)��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G@ϔ��ph!G��Ù���<ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�
mouseParam��editorCode.editorMousePivot��MousePivotParams���)��}�(j�  h)��}�(h G        h!G        ub�begin�h)��}�(h G@
��k]*Th!G���B�gub�end�h)��}�(h G@
��k]*Th!G����=�i@ub�dPivot�h)��}�(h G@
��k]*Th!G����=�i@ub�dEnd�h)��}�(h G        h!G�ѳf��Pub�dA�hA)��}�(hDG��s	6�hEG��.(�s�hFG?�����ub�dS�G?�Pu��ﴌangleOffset�G���bƠ��length�G@^@��hub�mode�K�active���obj�j�  ub�newObj�j   �
startPoint�h)��}�(h G?�4�H*��h!G?�V��hubj�  h)��}�(h G        h!G        ubj�  K�	processed���oldObjectAnchor�h)��}�(h G������?0h!G��g���ub�oldObjectAngle�hA)��}�(hDG        hEG        hFG?�      ub�oldObjectScale�G?�      ubj�  )��}�(j�  j`  hj�  j�  j   ubj�  )��}�(h,j�  j�  j�  j�  h)��}�(h G@
��k]*Th!G���B�gubj�  h)��}�(h G        h!G        ubj�  Kj�  �j�  h)��}�(h G@ϔ��ph!G��Ù���<ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(j�  j`  hhj�  j�  ubj�  )��}�(j�  j`  hj"  j�  hubj�  )��}�(j�  j`  hhj�  j   ubj�  )��}�(j�  j  j�  �j�  G        j�  G@i      ubj�  )��}�(j�  j`  hjF  j�  j\  ubj�  )��}�(jv  jD  j�  G@o@     j�  G@i      ubj�  )��}�(j�  j`  hj^  j�  jD  ubj�  )��}�(jv  j\  j�  G@o@     j�  G@i      ubjq  �ComCreateMapping���)��}�(j�  j`  hh�mapping�j(  �prevMapping�jt  ubjq  �ComSetMappingFromSelection���)��}�(j�  j(  �	selection�h�	Selection���)��}�(�start�h)��}�(h G@d�c�?c�h!G@M㻻���ubj�  h)��}�(h G@e������h!G@I�a�ubj�  �ub�	oldOffset�jO  �oldSize�jN  ubj�  )��}�(h,j�  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G?�D���>h!G?Ȇ`�P�ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?��mѤ\ubj�  j�  )��}�(j�  h)��}�(h G?�J�+x|h!G?��R�Youbj�  h)��}�(h G?�\�r<7h!G?�Ow֧�lubj�  h)��}�(h G?�V1����h!G?������ubj�  h)��}�(h G�Ϥ�.�m�h!G?��Z�ǝ�ubj�  h)��}�(h G���XN�+�h!G?�|�4�%�ubj�  hA)��}�(hDG���(�k�hhEG����x�hFG?�i-�i�ubj�  G@�o���j�  G� �k��bj�  G?�/RAubj�  Kj�  �j�  j(  ubj�  j(  j�  h)��}�(h G?�@h��&h!G?�oF]��ubj�  h)��}�(h G        h!G        ubj�  Kj�  �j�  h)��}�(h G        h!G        ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(j�  j(  j�  j�  j�  jO  j�  jN  ubjq  �ComSetPivot���)��}�(j�  jb  �newWorld�h)��}�(h G?�ۂ�Wz�h!G?՜�5�E�ub�oldWorld�h)��}�(h G        h!G        ububj�  )��}�(h,j   j�  j(  j�  h)��}�(h G?�>��h!G?��J���ubj�  h)��}�(h G?�J�+x|h!G?��R�Youbj�  Kj�  �j�  h)��}�(h G        h!G        ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�c&�+�cubj�  )��}�(j�  j(  j�  j�  j�  jO  j�  jN  ubj�  )��}�(h,j   j�  j(  j�  h)��}�(h G?��'�h!G?�Zx�3�ubj�  h)��}�(h G?�J�+x|h!G?��R�Youbj�  Kj�  �j�  h)��}�(h G?���ڔSDh!G?�����ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?���h:#ubj�  )��}�(j�  j(  j�  j�  j�  jO  j�  jN  ubj�  )��}�(h,j   j�  j(  j�  h)��}�(h G?�\�r<7h!G?�Ow֧�lubj�  h)��}�(h G?�J�+x|h!G?��R�Youbj�  Kj�  �j�  h)��}�(h G?�D���>h!G?Ȇ`�P�ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?��mѤ\ubj�  )��}�(j�  j(  j�  j�  j�  jO  j�  jN  ube�version��0.0.2�u.