��Y^      }�(�database��editorCode.database��Database���)��}�(�bodies�]�(�$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��	MainFrame��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G?�c���xh!G?�3�nFubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�>U��h!G?��֞?f<ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]��%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�c���xh!G?�3�nFububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�>U��h!G?��֞?f<ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1��
elasticity�G        �friction�G?�      �isSensor���shapeFilterGroup�K �shapeFilterCategory������ �shapeFilterMask������ �type��Polygon��internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G���sq3�8h!G?�L���ubh"h)��}�(h G���sq3�8h!G?�L���ububh)��}�(hh)��}�(h G��q q1��h!G?�0N䟠�ubh"h)��}�(h G��q q1��h!G?�0N䟠�ububh)��}�(hh)��}�(h G?궬���h!G?�~A��ubh"h)��}�(h G?궬���h!G?�~A��ububh)��}�(hh)��}�(h G?�����%�h!G?�@��*hubh"h)��}�(h G?�����%�h!G?�@��*hububh)��}�(hh)��}�(h G?���M�h!G?�ت�HV@ubh"h)��}�(h G?���M�h!G?�ت�HV@ububh)��}�(hh)��}�(h G��#�p�Hh!G?�&KɅvPubh"h)��}�(h G��#�p�Hh!G?�&KɅvPubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G?آ|�?bh!G?�HRS�ub�user�h)��}�(h G        h!G        ubh"h)��}�(h G?آ|�?bh!G?�HRS�ub�userDefined��ub�area�G?�4 �=��density�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h��ub�mass�h�)��}�(h�G?�      h�G@>      h"G@>      h��ub�moment�h�)��}�(h�G@#�zas{jh�G        h"G@#�zas{jh��ubububahl�Dynamic�h��+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G?آ|�?bh!G?�HRS�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?آ|�?bh!G?�HRS�ubh��ubh�G?�4 �=��h�h�)��}�(h�G@3�Dz�`h�G        h"G        h��ubh�h�)��}�(h�G@>      h�G        h"G@>      h��ubh�h�)��}�(h�G@#�zas{jh�G        h"G@#�zas{jh��ubububh)��}�(h�Wheel�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���ҶFfh!G����@&Vububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�rk#�#8h!G?�rk#�#8ubububh,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G�       h8G���ҶFfh9G        h:G?�rk#�#9h;G����@&Vubh<h)��}�(h G���ҶFfh!G����@&Vubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�rk#�#9ubhH]�hJ�Circle���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���ҶFfh!G����@&Vububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�rk#�#8h!G?�rk#�#8ubububh,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G�       h8G���ҶFfh9G        h:G?�rk#�#9h;G����@&Vubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE�hfG        hgG?�      hh�hiK hj����� hk����� hl�Circle�hnho�
CircleSpec���)��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G���ҶFfh!G����@&Vububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj  �radiusVector�h)��}�(h G        h!G        ubh�h�CircleRadius���)��}�(h"G?�rk#�#9�base�G?�      ub�	drawLines�K ubh�h��CirclePhysics���)��}�(h�h�)��}�(h�h)��}�(h G���ҶFfh!G����@&Vubh�h)��}�(h G        h!G        ubh"h)��}�(h G���ҶFfh!G����@&Vubh��ubh�G?��Q4�4h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@$      h"G@$      h��ubh�h�)��}�(h�G@	Kx�� h�G        h"G@	Kx�� h��ubububahlh�h�h�)��}�(h�h�)��}�(h�h)��}�(h G���ҶFfh!G����@&Vubh�h)��}�(h G        h!G        ubh"h)��}�(h G���ҶFfh!G����@&Vubh��ubh�G?��Q4�4h�h�)��}�(h�G@"h
���h�G        h"G        h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubh�h�)��}�(h�G@	Kx�� h�G        h"G@	Kx�� h��ubububh)��}�(h�Wheel_1�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?����HP�h!G���|䥄ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�rk#�#8h!G?�rk#�#8ubububh,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G�       h8G?����HP�h9G        h:G?�rk#�#9h;G���|䥄ubh<h)��}�(h G?����HP�h!G���|䥄ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�rk#�#9ubhH]�h�)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?����HP�h!G���|䥄ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�rk#�#8h!G?�rk#�#8ubububh,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G�       h8G?����HP�h9G        h:G?�rk#�#9h;G���|䥄ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfG        hgG?�      hh�hiK hj����� hk����� hl�Circle�hnj  )��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G?����HP�h!G���|䥄ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj}  j  h)��}�(h G        h!G        ubh�j  )��}�(h"G?�rk#�#9j"  G?�      ubj#  K ubh�j%  )��}�(h�h�)��}�(h�h)��}�(h G?����HP�h!G���|䥄ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?����HP�h!G���|䥄ubh��ubh�G?��Q4�4h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@$      h"G@$      h��ubh�h�)��}�(h�G@	Kx�� h�G        h"G@	Kx�� h��ubububahl�Dynamic�h�h�)��}�(h�h�)��}�(h�h)��}�(h G?����HP�h!G���|䥄ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?����HP�h!G���|䥄ubh��ubh�G?��Q4�4h�h�)��}�(h�G@"h
���h�G        h"G        h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubh�h�)��}�(h�G@	Kx�� h�G        h"G@	Kx�� h��ububube�	shapeList�]�(h�hMj`  e�constraints�]�(�/editorCode.constraintInternals.editorConstraint��DampedSpring���)��}�(h�CNSTRNT�hl�Damped Spring��bodyA�h�bodyB�hԌselfCollide���maxForce�G�      �maxBias�G�      �	errorBias�G?]q5�NZ�
restLength�G        �	stiffness�G@@     �damping�G@D      �anchorA�h�OffsetPoint���)��}�(�offset�h)��}�(h G�����
h!G�����3{Bubhh)��}�(h G�����
h!G�����3{Bubh"h)��}�(h G��ֿ�A8|h!G��N��
QKubub�anchorB�j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���ҶFfh!G����@&Vubububj�  �GrooveJoint���)��}�(h�	CNSTRNT_1�hl�Groove�j�  hj�  h�j�  �j�  G�      j�  G�      j�  G?]q5�NZ�grooveA�j�  )��}�(j�  h)��}�(h G�����h!G��/�ò��ubhh)��}�(h G�����h!G��/�ò��ubh"h)��}�(h G���Z�7gvh!G?��BT�K`ubub�grooveB�j�  )��}�(j�  h)��}�(h G��� �th!G��b��'O%ubhh)��}�(h G��� �th!G��b��'O%ubh"h)��}�(h G����qaPh!G��W��%.ububj�  j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���ҶFfh!G����@&Vubububj�  )��}�(h�	CNSTRNT_2�hl�Damped Spring�j�  hj�  jF  j�  �j�  G�      j�  G�      j�  G?]q5�NZj�  G        j�  G@@     j�  G@D      j�  j�  )��}�(j�  h)��}�(h G?�.F��Hdh!G���n����ubhh)��}�(h G?�.F��Hdh!G���n����ubh"h)��}�(h G?�V��i�h!G��Zʱj}�ububj�  j�  )��}�(j�  h)��}�(h G�k<�B��h!G?u��Xl��ubhh)��}�(h G�e���J� h!G?q?X#  ubh"h)��}�(h G?��vh+5h!G���Dz���ubububj�  )��}�(h�	CNSTRNT_3�hl�Groove�j�  hj�  jF  j�  �j�  G�      j�  G�      j�  G?]q5�NZj�  j�  )��}�(j�  h)��}�(h G?��a��/�h!G���pqG�ubhh)��}�(h G?��a��/�h!G���pqG�ubh"h)��}�(h G?�� ڳ�ph!G?��L�ububj�  j�  )��}�(j�  h)��}�(h G?�]�u���h!G������Mubhh)��}�(h G?�]�u���h!G������Mubh"h)��}�(h G?�������h!G���f�Vububj�  j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G?����HP�h!G���|䥄ububube�mappings�]�(�editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�      h!G��      ubh"h)��}�(h G�      h!G��      ububh)��}�(hh)��}�(h G@      h!G��      ubh"h)��}�(h G@      h!G��      ububh)��}�(hh)��}�(h G�      h!G?�      ubh"h)��}�(h G�      h!G?�      ububh)��}�(hh)��}�(h G@      h!G?�      ubh"h)��}�(h G@      h!G?�      ubube�textureSize�]�(K�K`e�anchor�]�(G@X      G@H      e�mappingSize�]�(K�K`e�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@[O����h!G@Q�����ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububj+  )��}�(h�MAP:1�j/  Kj0  h�h,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G        h8G���ҶFfh9G        h:G?�rk#�#9h;G����@&Vubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj9  ]�(h)��}�(hh)��}�(h G��      h!G        ubh"h)��}�(h G�H$�h!G����@&Vububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G���$f��h!G����@&Vububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G�H$�h!G���A��R�ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G���$f��h!G���A��R�ububejS  ]�(K@K@ejU  ]�(G@@      G@@      ejW  ]�(K@K ejY  ]�(K K ej[  ]�(h)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubjg  h)��}�(hh)��}�(h G        h!G?�      ubh"h)��}�(h G���ҶFfh!G��0�f��ubububj+  )��}�(h�	MAP:1_1:2�j/  Kj0  h�h,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G        h8G���ҶFfh9G        h:G?�rk#�#9h;G����@&Vubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj9  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G�H$�h!G���;���ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G���$f��h!G���;���ububh)��}�(hh)��}�(h G��      h!G        ubh"h)��}�(h G�H$�h!G����@&Vububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G���$f��h!G����@&VububejS  ]�(K@K@ejU  ]�(G@@      G@@      ejW  ]�(K@K ejY  ]�(K K ej[  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubjg  h)��}�(hh)��}�(h G        h!G��      ubh"h)��}�(h G���ҶFfh!G��Q��/�$ubububj+  )��}�(h�MAP:1:1�j/  Kj0  jF  h,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G        h8G?����HP�h9G        h:G?�rk#�#9h;G���|䥄ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj9  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?�үWh��h!G�����ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@"�=��h!G�����ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G?�үWh��h!G�ԭ7�O�ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G@"�=��h!G�ԭ7�O�ububejS  ]�(K@K@ejU  ]�(G@@      G@@      ejW  ]�(K@K"ejY  ]�(K Kej[  ]�(h)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubjg  h)��}�(hh)��}�(h G        h!G?�      ubh"h)��}�(h G?����HP�h!G���d���ubububj+  )��}�(h�MAP:1_1:2:2�j/  Kj0  jF  h,h.)��}�(h1h3)��}�(h6G?�rk#�#9h7G        h8G?����HP�h9G        h:G?�rk#�#9h;G���|䥄ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj9  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?�үWh��h!G�����7 ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@"�=��h!G�����7 ububh)��}�(hh)��}�(h G��      h!G        ubh"h)��}�(h G?�үWh��h!G���|䥄ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G@"�=��h!G���|䥄ububejS  ]�(K@K@ejU  ]�(G@@      G@@      ejW  ]�(K@K ejY  ]�(K K ej[  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubjg  h)��}�(hh)��}�(h G        h!G��      ubh"h)��}�(h G?����HP�h!G��AE�nRubububeub�textureSizes�]�(K�K`��K@K@��K@K@��K K ��jW  jW  jW  jW  jW  jW  jW  jW  jW  jW  jW  jW  e�texturePaths�]�(�data\textures\truck.png��data\textures\wheel1.png��data\textures\wheel2.png�� �j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�hԌcurrentShape�h��currentConstraint�j�  �currentMapping�j�  �currentMappingChannel�Khh)��}�(hhj�  j�  j�  j�  j'  j(  ububhjt  �object�h�prevCurrent�Nubjf  )��}�(ji  jm  hjt  jv  h�jw  hubjd  �ComSetBodyAsCurrent���)��}�(ji  jm  h�BODY_1��prev�h�ubjd  �ComRenameBody���)��}�(j0  h�hjt  �newName�h֌oldName�j~  ubj{  )��}�(ji  jm  h�BODY�j  h�ubjd  �ComStartTransform���)��}�(h,�editorCode.editorViewTransform��ContinuousTransform���)��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G����>��h!G�������ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�
mouseParam��editorCode.editorMousePivot��MousePivotParams���)��}�(�pivot�h)��}�(h G���xϦCh!G������`�ub�begin�h)��}�(h G��1o��
h!G?���MǼub�end�h)��}�(h G�	�l'}�&h!G?��&Őub�dPivot�h)��}�(h G��_T�4h!G?��lL�9�ub�dEnd�h)��}�(h G?̬T��@h!G��1��,�ub�dA�hA)��}�(hDG?��r|��hEG?�١�ZJhFG?���`�|�ub�dS�G?�rk#�#9�angleOffset�G@��|��t�length�G@�^1Lub�mode�K�active���obj�h�ub�newObj�h�
startPoint�h)��}�(h G@����h!G?�$�I$�Hubj�  h)��}�(h K h!K ubj�  K�	processed���oldObjectAnchor�h)��}�(h G        h!G        ub�oldObjectAngle�hA)��}�(hDG        hEG        hFG?�      ub�oldObjectScale�G?�      ubj�  )��}�(h,j�  j�  hj�  h)��}�(h G@����h!G?�$�I$�Hubj�  h)��}�(h K h!K ubj�  K j�  �j�  h)��}�(h G        h!G        ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(h,j�  j�  hj�  h)��}�(h G@����h!G?�$�I$�Hubj�  h)��}�(h K h!K ubj�  Kj�  �j�  h)��}�(h G        h!G        ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(j0  hhjt  j�  hj�  j�  ubj{  )��}�(ji  jm  hh�j  hubjd  �ComLoadTexture���)��}�(hjt  �newPath�jZ  �destChannel�K �newSize�jT  �oldPath�j]  �oldSize�jW  ubj�  )��}�(hjt  j�  j[  j�  Kj�  jU  j�  j]  j�  jW  ubjd  �ComCreateMapping���)��}�(ji  jm  hjt  �mapping�j,  �prevMapping�Nubj�  )��}�(ji  jm  hjt  j�  jn  j�  Nubj�  )��}�(ji  jm  hjt  j�  j+  )��}�(h�MAP:1_1�j/  Kj0  Nh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj9  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G        h!G        ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G        h!G        ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G        h!G        ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G        h!G        ububejS  ]�(K@K@ejU  ]�(G@@      G@@      ejW  ]�(K@K@ejY  ]�(K K ej[  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G        h!G        ubjg  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububj�  jn  ubjd  �ComDeleteMapping���)��}�(ji  jm  hjt  j�  j�  �index�K�current��ubj{  )��}�(ji  jm  hhj  h�ubj{  )��}�(ji  jm  hh�j  hubj{  )��}�(ji  jm  hh�j  h�ubjd  �ComAddNewShape���)��}�(ji  jm  hjt  �shape�h��	prevShape�Nj0  h�ubj{  )��}�(ji  jm  hhj  h�ubj9  )��}�(ji  jm  hjt  j<  hMj=  Nj0  hubjd  �ComNewShapeAddPoint���)��}�(j<  hM�point�hvubjC  )��}�(j<  hMjF  h|ubjC  )��}�(j<  hMjF  h�ubjC  )��}�(j<  hMjF  h�ubjC  )��}�(j<  hMjF  h�ubjC  )��}�(j<  hMjF  h�ubjd  �ComSetUserParam���)��}�(�param�h��oldUserFlag���
oldUserVal�G        �value�G@>      ubjd  �ComSelectNextBody���)��}�(ji  jm  �oldBody�h�oldShape�hM�newBody�hԌnewShape�h��executed��ubjR  )��}�(jU  j2  jV  �jW  G        jX  G@$      ubj{  )��}�(ji  jm  hh�j  h�ubj�  )��}�(h,j�  j�  h�j�  h)��}�(h G?��<0��|h!G?��̨�1�ubj�  h)��}�(h K h!K ubj�  Kj�  �j�  h)��}�(h G        h!G        ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubj�  )��}�(h,j�  j�  h�j�  h)��}�(h G��$�aռh!G�� `��8ubj�  h)��}�(h K h!K ubj�  Kj�  �j�  h)��}�(h G��9ʹX�h!G��Rg~`ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubjd  �ComSetPivot���)��}�(j�  h)��}�(h G���xϦCh!G������`�ub�newWorld�h)��}�(h G���xϦCh!G������`�ub�oldWorld�h)��}�(h K h!K ububj�  )��}�(h,j�  j�  h�j�  h)��}�(h G��7˖@h!G?��+;�� ubj�  h)��}�(h G���xϦCh!G������`�ubj�  Kj�  �j�  h)��}�(h G��k2w��h!G�О ���ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubjd  �ComSetMappingFromSelection���)��}�(j�  jn  �	selection�h�	Selection���)��}�(�start�h)��}�(h G��X-@�h!G@?�{1?1rubj�  h)��}�(h G@P6��ߋh!G�+#����ubj�  �ub�	oldOffset�j�  j�  j�  ubj�  )��}�(j�  jn  j�  j�  j�  j�  j�  j�  ubj�  )��}�(hjt  j�  j\  j�  Kj�  jV  j�  j]  j�  jW  ubj�  )��}�(ji  jm  hjt  j�  j�  j�  Nubj�  )��}�(j�  j�  j�  j�  j�  j�  j�  j�  ubj�  )��}�(h,j�  j�  h�j�  h)��}�(h G��1o��
h!G?���MǼubj�  h)��}�(h G���xϦCh!G������`�ubj�  Kj�  �j�  h)��}�(h G����>��h!G�������ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�      ubjd  �ComAddConstraint���)��}�(hjt  ji  jm  jv  j�  jw  Nubjd  �ComConstraintSetNewBodyA���)��}�(�entity�j�  j_  hj]  Nubj�  )��}�(j�  j�  j_  h�j]  hubj�  )��}�(j�  j�  j_  hj]  h�ubjd  �ComConstraintSetNewBodyB���)��}�(j�  j�  j_  h�j]  Nubjd  �ComSetAnchorAFromCoords���)��}�(j�  j�  �	newXValue�G��ſ��	newYValue�G��� �㭌	oldXValue�G        �	oldYValue�G        ubj�  )��}�(j�  j�  j�  G����#��j�  G��!�P�B�j�  G��ſ�j�  G��� ��ubj�  )��}�(j�  j�  j�  G����#��j�  G��!�P�B�j�  G����#��j�  G��!�P�B�ubj�  )��}�(j�  j�  j�  G��#�A!j�  G��%0��.j�  G����#��j�  G��!�P�B�ubj�  )��}�(j�  j�  j�  G��#�A!j�  G��%0��.j�  G��#�A!j�  G��%0��.ubj�  )��}�(j�  j�  j�  G����#��j�  G��)B#�~j�  G��#�A!j�  G��%0��.ubj�  )��}�(j�  j�  j�  G���k�j�  G��CL*X1�j�  G����#��j�  G��)B#�~ubj�  )��}�(j�  j�  j�  G��@�9Ɛj�  G��CY"�`uj�  G���k�j�  G��CL*X1�ubj�  )��}�(j�  j�  j�  G��x+�#Mj�  G��CY"�`uj�  G��@�9Ɛj�  G��CY"�`uubj�  )��}�(j�  j�  j�  G� :�9�j�  G��CY"�`uj�  G��x+�#Mj�  G��CY"�`uubj�  )��}�(j�  j�  j�  G��x+�#Mj�  G��C��^�j�  G� :�9�j�  G��CY"�`uubj�  )��}�(j�  j�  j�  G��q9��j�  G����4�j�  G��x+�#Mj�  G��C��^�ubj�  )��}�(j�  j�  j�  G������tj�  G����4�j�  G��q9��j�  G����4�ubj�  )��}�(j�  j�  j�  G������j�  G����W��5j�  G������tj�  G����4�ubj�  )��}�(j�  j�  j�  G����͚$j�  G����W��5j�  G������j�  G����W��5ubj�  )��}�(j�  j�  j�  G��cg�S�j�  G����W��5j�  G����͚$j�  G����W��5ubj�  )��}�(j�  j�  j�  G��@�9Ɛj�  G�����3{Bj�  G��cg�S�j�  G����W��5ubj�  )��}�(j�  j�  j�  G�����
j�  G�����3{Bj�  G��@�9Ɛj�  G�����3{Bubjd  �ComSetRestLength���)��}�(j�  j�  �newValue�G        �oldValue�G?�      ubjd  �ComSetDamping���)��}�(j�  j�  j�  G@D      j�  G?�      ubjd  �ComSetStiffness���)��}�(j�  j�  j�  G@@     j�  G?�      ubj�  )��}�(hjt  ji  jm  jv  j�  jw  j�  ubj�  )��}�(j�  j�  j_  hj]  Nubj�  )��}�(j�  j�  j_  h�j]  Nubjd  �ComSetGrooveBFromCoords���)��}�(j�  j�  j�  G��� �tj�  G��b��'O%j�  G        j�  G        ubjd  �ComSetGrooveAFromCoords���)��}�(j�  j�  j�  G�����j�  G��/�ò��j�  G        j�  G        ubj{  )��}�(ji  jl  )��}�(jo  h�jp  h�jq  j�  jr  jn  js  Khh)��}�(hhj�  j�  j�  j�  j'  j(  ububhh�j  h�ubjd  �ComBodyClone���)��}�(�baseBody�h�hj  j_  jF  �preRun��hH]�j`  a�newConstraintsA�]��newConstraintsB�]�(j�  j  e�newMappings�]�(j�  j  eubj�  )��}�(h,j�  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G?�,]zh!G����� ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�rk#�#9ubj�  j�  )��}�(j�  h)��}�(h G?���C�Vhh!G���4��Šubj�  h)��}�(h G?�踲{�(h!G���&g��&ubj�  h)��}�(h G@K���\h!G��B��ubj�  h)��}�(h G?��XRW��h!G?�1^Q�ubj�  h)��}�(h G?�N��H�h!G?ޔvJ��pubj�  hA)��}�(hDG����shEG��n�R�-hFG������Y[ubj�  G?�o^�_?j�  G�����j�  G?�oIHgubj�  Kj�  �j�  jF  ubj�  jF  j�  h)��}�(h G�������h!G?�k
|���ubj�  h)��}�(h K h!K ubj�  Kj�  �j�  h)��}�(h G���ҶFfh!G����@&Vubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�rk#�#9ubj{  )��}�(j�  h)��}�(h G?���C�Vhh!G���4��Šubj�  h)��}�(h G?���C�Vhh!G���4��Šubj�  h)��}�(h K h!K ububj�  )��}�(h,j  j�  jF  j�  h)��}�(h G?�踲{�(h!G���&g��&ubj�  h)��}�(h G?���C�Vhh!G���4��Šubj�  Kj�  �j�  h)��}�(h G?�,]zh!G����� ubj�  hA)��}�(hDG        hEG        hFG?�      ubj�  G?�rk#�#9ubjZ  )��}�(ji  j
  j]  jF  j^  j`  j_  hj`  hMja  �ubjZ  )��}�(ji  j
  j]  hj^  hMj_  h�j`  h�ja  �ubj�  )��}�(j�  jn  j�  j�  )��}�(j�  h)��}�(h G�����h!G@P�viik�ubj�  h)��}�(h G@P�_�e�h!G@@��s3 ubj�  �ubj�  j�  j�  j�  ubjd  �ComSetConstraintAsCurrent���)��}�(ji  j
  hj  j  j�  ubj\  )��}�(ji  j
  hj�  j  j  ubjd  �ComSetRestLengthFromCoords���)��}�(j�  G@�l�{�j�  j�  j�  G        ubjb  )��}�(j�  G@����j�  j�  j�  G@�l�{�ubjb  )��}�(j�  G@�:&j�  j�  j�  G@����ubjb  )��}�(j�  G@����j�  j�  j�  G@�:&ubjb  )��}�(j�  G@s��Xj�  j�  j�  G@����ubjb  )��}�(j�  G@�	��Aj�  j�  j�  G@s��Xubjb  )��}�(j�  G@�<��kj�  j�  j�  G@�	��Aubjb  )��}�(j�  G@��ڎAj�  j�  j�  G@�<��kubjb  )��}�(j�  G@r�j�  j�  j�  G@��ڎAubjb  )��}�(j�  G@���ej�  j�  j�  G@r�ubjb  )��}�(j�  G@��X>oj�  j�  j�  G@���eubjb  )��}�(j�  G@��,=��j�  j�  j�  G@��X>oubjb  )��}�(j�  G@��,=��j�  j�  j�  G@��,=��ubjb  )��}�(j�  G@���I�j�  j�  j�  G@��,=��ubjb  )��}�(j�  G@��f'��j�  j�  j�  G@���I�ubjd  �ComSetAnchorBFromCoords���)��}�(j�  j�  j�  G?8�]2j�  G?��4�*t�j�  G        j�  G        ubj�  )��}�(j�  j�  j�  G?8�]2j�  G?�����Aj�  G?8�]2j�  G?��4�*t�ubj�  )��}�(j�  j�  j�  G�k<�B��j�  G?u��Xl��j�  G?8�]2j�  G?�����Aubj�  )��}�(j�  j�  j�  G?�Rk!��j�  G���z�JA�j�  G�����
j�  G�����3{Bubj�  )��}�(j�  j�  j�  G?�^wOs��j�  G��ȇ ��j�  G?�Rk!��j�  G���z�JA�ubj�  )��}�(j�  j�  j�  G?�.F��Hdj�  G���n����j�  G?�^wOs��j�  G��ȇ ��ubj�  )��}�(j�  j�  j�  G        j�  G@��f'��ubj�  )��}�(j�  jn  j�  jU  j�  j�  j�  j�  ubj�  )��}�(j�  jn  j�  jU  j�  j�  j�  j�  ubj�  )��}�(j�  jn  j�  jU  j�  j�  j�  j�  ubj\  )��}�(ji  jl  )��}�(jo  jF  jp  j`  jq  j�  jr  j  js  Khhubhj  j  j  ubj\  )��}�(ji  j�  hj�  j  j  ubj\  )��}�(ji  j�  hj�  j  j�  ubj\  )��}�(ji  j�  hj  j  j�  ubj  )��}�(j�  j  j�  G?�]�u���j�  G������Mj�  G��� �tj�  G��b��'O%ubj  )��}�(j�  j  j�  G?�J�b��j�  G���ԘvMnj�  G�����j�  G��/�ò��ubj  )��}�(j�  j  j�  G?��a��/�j�  G���pqG�j�  G?�J�b��j�  G���ԘvMnubj\  )��}�(ji  j�  hj  j  j  ubj\  )��}�(ji  j�  hj  j  j  ubj\  )��}�(ji  j�  hj�  j  j  ubj\  )��}�(ji  j�  hj�  j  j�  ubj\  )��}�(ji  j�  hj�  j  j�  ube�version��0.0.2�u.