��R      }�(�database��editorCode.database��Database���)��}�(�bodies�]��$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��BODY��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G        h!G        ubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G        h!G        ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]��%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�333330h!G?�:��<ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�PuPuh!G?�PuPuubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��type�hK�internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G��A�A�h!G��A�A� ubh"h)��}�(h G��A�A�h!G��A�A� ububh)��}�(hh)��}�(h G��333334h!G?�������ubh"h)��}�(h G��333334h!G?�������ububh)��}�(hh)��}�(h G��ffffffh!G?䯊����ubh"h)��}�(h G��ffffffh!G?䯊����ububh)��}�(hh)��}�(h G�è:��:�h!G?�PuPuubh"h)��}�(h G�è:��:�h!G?�PuPuububh)��}�(hh)��}�(h G?ϊ�����h!G?�:��:�ubh"h)��}�(h G?ϊ�����h!G?�:��:�ububh)��}�(hh)��}�(h G?��_�_h!G?�:��:�ubh"h)��}�(h G?��_�_h!G?�:��:�ububh)��}�(hh)��}�(h G?噙����h!G?�����ubh"h)��}�(h G?噙����h!G?�����ububh)��}�(hh)��}�(h G?惨:��:h!G?�W�|W�|ubh"h)��}�(h G?惨:��:h!G?�W�|W�|ububh)��}�(hh)��}�(h G?�������h!G��A�A�ubh"h)��}�(h G?�������h!G��A�A�ububh)��}�(hh)��}�(h G?��A�Bh!G���_�^ubh"h)��}�(h G?��A�Bh!G���_�^ububh)��}�(hh)��}�(h G?�A�A�h!G��_�_�ubh"h)��}�(h G?�A�A�h!G��_�_�ububh)��}�(hh)��}�(h G��I$�I$�h!G��ffffffubh"h)��}�(h G��I$�I$�h!G��ffffffububh)��}�(hh)��}�(h G��PuPuh!G�ொ����ubh"h)��}�(h G��PuPuh!G�ொ����ububh)��}�(hh)��}�(h G���+�,h!G�د�����ubh"h)��}�(h G���+�,h!G�د�����ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G?�����M3h!G?��OA��ub�user�h)��}�(h G        h!G        ubh"h)��}�(h G?�����M3h!G?��OA��ub�userDefined��ub�area�G?���v�یdensity�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h܉ub�mass�h�)��}�(h�G?�      h�G        h"G?���v��h܉ub�moment�h�)��}�(h�G?ۚY!�`h�G        h"G?ۚY!�`h܉ubububahf�Dynamic�hɌ+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G        h!G        ubh�h)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubh܉ubh�G?�      h�h�)��}�(h�G?�      h�G        h"G?�      h܉ubh�h�)��}�(h�G?�      h�G        h"G?�      h܉ubh�h�)��}�(h�G?�      h�G        h"G?�      h܉ubububa�	shapeList�]�hMa�constraints�]��mappings�]�ub�textureSizes�]�(K K ��j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  e�texturePaths�]�(� �j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  e�queueProcessed��collections��deque���)Kd��R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�h�currentShape�hM�currentConstraint�N�currentMapping�N�currentMappingChannel�K hhubhh�object�h�prevCurrent�Nubj  �ComAddNewShape���)��}�(j  j  hh�shape�hM�	prevShape�N�body�hubj  �ComNewShapeAddPoint���)��}�(j%  hM�point�houbj)  )��}�(j%  hMj,  huubj)  )��}�(j%  hMj,  h{ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubj)  )��}�(j%  hMj,  h�ubeu.