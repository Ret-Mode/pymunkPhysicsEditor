���k      }�(�database��editorCode.database��Database���)��}�(�bodies�]�(�$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��Main��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G?����K h!G?�c�1�ubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@x���yh!G?�+����\ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]��%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?����K h!G?�c�1�ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@x���yh!G?�+����\ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��type��Polygon��internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G@�����h!G��A4e�ubh"h)��}�(h G@�����h!G��A4e�ububh)��}�(hh)��}�(h G?��;7Th!G���'�ubh"h)��}�(h G?��;7Th!G���'�ububh)��}�(hh)��}�(h G��3c%W4�h!G���v��E�ubh"h)��}�(h G��3c%W4�h!G���v��E�ububh)��}�(hh)��}�(h G���G��՜h!G���'�ubh"h)��}�(h G���G��՜h!G���'�ububh)��}�(hh)��}�(h G��I1j h!G���56�6Hubh"h)��}�(h G��I1j h!G���56�6Hububh)��}�(hh)��}�(h G�c�E� .h!G?Εد]O ubh"h)��}�(h G�c�E� .h!G?Εد]O ububh)��}�(hh)��}�(h G�����Mh!G?���ީ��ubh"h)��}�(h G�����Mh!G?���ީ��ububh)��}�(hh)��}�(h G��fm��)�h!G?���[jlubh"h)��}�(h G��fm��)�h!G?���[jlububh)��}�(hh)��}�(h G��O����h!G?��!�%(�ubh"h)��}�(h G��O����h!G?��!�%(�ububh)��}�(hh)��}�(h G?ԃB�h!G?��G���ubh"h)��}�(h G?ԃB�h!G?��G���ububh)��}�(hh)��}�(h G?�x_4z�h!G?�Q(�Wz�ubh"h)��}�(h G?�x_4z�h!G?�Q(�Wz�ububh)��}�(hh)��}�(h G?��s���h!G?�$�$�� ubh"h)��}�(h G?��s���h!G?�$�$�� ububh)��}�(hh)��}�(h G@VCު�h!G?�1;׏ubh"h)��}�(h G@VCު�h!G?�1;׏ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G��	,�̷�h!G?�ɱ�C�?ub�user�h)��}�(h G        h!G        ubh"h)��}�(h G��	,�̷�h!G?�ɱ�C�?ub�userDefined��ub�area�G@q)�h��density�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h׉ub�mass�h�)��}�(h�G?�      h�G        h"G@q)�h�h׉ub�moment�h�)��}�(h�G@0��6P��h�G        h"G@0��6P��h׉ubububahf�Dynamic�hČ+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G��	,�̷�h!G?�ɱ�C�?ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��	,�̷�h!G?�ɱ�C�?ubh׉ubh�G@q)�h�h�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G@q)�h�h�G        h"G@q)�h�h׉ubh�h�)��}�(h�G@0��6P��h�G        h"G@0��6P��h׉ubububh)��}�(h�WHeelL�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G��,��h!G���T��~�ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G��,��h9G        h:G?�      h;G���T��~�ubh<h)��}�(h G��,��h!G���T��~�ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�hJ�Circle���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G��,��h!G���T��~�ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G��,��h9G        h:G?�      h;G���T��~�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1�hf�Circle�hhhi�
CircleSpec���)��}�(hn]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G��,��h!G���T��~�ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj3  �radiusVector�h)��}�(h G        h!G        ubh�h�CircleRadius���)��}�(h"G?�      �base�G?�      ub�	drawLines�K ubh�hŌCirclePhysics���)��}�(h�h�)��}�(h�h)��}�(h G��,��h!G���T��~�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��,��h!G���T��~�ubh׉ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h׉ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h׉ubububahfh�h�h�)��}�(h�h�)��}�(h�h)��}�(h G��,��h!G���T��~�ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��,��h!G���T��~�ubh׉ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G@	!�TD-h�G        h"G@	!�TD-h׉ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h׉ubububh)��}�(h�WHeelR�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�U��Hih!G��Ƅ���ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G@�U��Hih9G        h:G?�      h;G��Ƅ���ubh<h)��}�(h G@�U��Hih!G��Ƅ���ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�j  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�U��Hih!G��Ƅ���ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G@�U��Hih9G        h:G?�      h;G��Ƅ���ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfj-  hhj/  )��}�(hn]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@�U��Hih!G��Ƅ���ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj�  j?  h)��}�(h G        h!G        ubh�jC  )��}�(h"G?�      jF  G?�      ubjG  K ubh�jI  )��}�(h�h�)��}�(h�h)��}�(h G@�U��Hih!G��Ƅ���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@�U��Hih!G��Ƅ���ubh׉ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G?�      h�G        h"G@	!�TD-h׉ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h׉ubububahfh�h�h�)��}�(h�h�)��}�(h�h)��}�(h G@�U��Hih!G��Ƅ���ubh�h)��}�(h G        h!G        ubh"h)��}�(h G@�U��Hih!G��Ƅ���ubh׉ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G@	!�TD-h�G        h"G@	!�TD-h׉ubh�h�)��}�(h�G?�!�TD-h�G        h"G?�!�TD-h׉ububube�	shapeList�]�(hMj  j�  e�constraints�]�(�/editorCode.constraintInternals.editorConstraint��GrooveJoint���)��}�(h�CNSTRNT�hf�Groove��bodyA�h�bodyB�h��collideBodies���	max_force�G?�      �grooveA�h�OffsetPoint���)��}�(�offset�h)��}�(h G��W��[Lh!G��W�$@ubhh)��}�(h G��W��[Lh!G��W�$@ubh"h)��}�(h G��`�G(h!G����8�Rpubub�grooveB�j�  )��}�(j�  h)��}�(h G��W��[Lh!G?�J�y��ubhh)��}�(h G��W��[Lh!G?�J�y��ubh"h)��}�(h G��`�G(h!G?�}>�`�(ubub�anchorB�j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G��,��h!G���T��~�ubububj�  )��}�(h�	CNSTRNT_1�hfj�  j�  hj�  jj  j�  �j�  G?�      j�  j�  )��}�(j�  h)��}�(h G@���Mh!G��6��>�4ubhh)��}�(h G@���Mh!G��6��>�4ubh"h)��}�(h G@�h�dh!G��:�=��Xububj�  j�  )��}�(j�  h)��}�(h G@	z:�!Ph!G?�rCaɐubhh)��}�(h G@	z:�!Ph!G?�rCaɐubh"h)��}�(h G@�q-T�h!G?꤆�2��ububj�  j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@�U��Hih!G��Ƅ���ubububj�  �DampedSpring���)��}�(h�	CNSTRNT_2�hf�Damped Spring�j�  hj�  h�j�  �j�  G?�      �
restLength�G        �	stiffness�G@@     �damping�G@4      �anchorA�j�  )��}�(j�  h)��}�(h G��i�8h!G�}��ubhh)��}�(h G��i�8h!G�}��ubh"h)��}�(h G��#5��h!G��u:����ububj�  j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G��,��h!G���T��~�ubububj  )��}�(h�	CNSTRNT_3�hfj  j�  hj�  jj  j�  �j�  G?�      j  G        j  G@@     j   G@4      j!  j�  )��}�(j�  h)��}�(h G@=� h!G��d첾\ubhh)��}�(h G@=� h!G��d첾\ubh"h)��}�(h G@�3�93`h!G����u��Lububj�  j�  )��}�(j�  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G@�U��Hih!G��Ƅ���ububube�mappings�]�(�editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�      h!G��      ubh"h)��}�(h G�      h!G��      ububh)��}�(hh)��}�(h G@      h!G��      ubh"h)��}�(h G@      h!G��      ububh)��}�(hh)��}�(h G�      h!G?�      ubh"h)��}�(h G�      h!G?�      ububh)��}�(hh)��}�(h G@      h!G?�      ubh"h)��}�(h G@      h!G?�      ubube�textureSize�]�(K�K`e�anchor�]�(G@X      G@H      e�mappingSize�]�(K�K`e�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@X      h!G@H      ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububjI  )��}�(h�MAP:1�jM  KjN  h�h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G��,��h9G        h:G?�      h;G���T��~�ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubjW  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G��,��h!G����N?Hububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G���Y=hh!G����N?Hububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G��,��h!G?�%V��ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G���Y=hh!G?�%V��ububejq  ]�(K@K@ejs  ]�(G@@      G@@      eju  ]�(K@K@ejw  ]�(K K ejy  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G��,��h!G���T��~�ubububjI  )��}�(h�MAP:1_1�jM  KjN  jj  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G@�U��Hih9G        h:G?�      h;G��Ƅ���ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubjW  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?������h!G��cB~��]ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@�U��Hih!G��cB~��]ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G?������h!G?�r�"�ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G@�U��Hih!G?�r�"�ububejq  ]�(K@K@ejs  ]�(G@@      G@@      eju  ]�(K@K@ejw  ]�(K K ejy  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G@�U��Hih!G��Ƅ���ubububeub�textureSizes�]�(K�K`��K@K@��K K ��j  j  j  j  j  j  j  j  j  j  j  j  j  e�texturePaths�]�(�data/textures/pinky.png��data/textures/wheel2.png�� �j  j  j  j  j  j  j  j  j  j  j  j  j  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�jj  �currentShape�j�  �currentConstraint�j�  �currentMapping�j�  �currentMappingChannel�Khh)��}�(hhj�  j�  j�  j�  jE  jF  ububhj  �object�h�prevCurrent�Nubj  )��}�(j  j  hj  j   h�j!  hubj  �ComStartTransform���)��}�(h,�editorCode.editorViewTransform��ContinuousTransform���)��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G@$��W�h!G���N�1�ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�
mouseParam��editorCode.editorMousePivot��MousePivotParams���)��}�(�pivot�h)��}�(h K h!K ub�begin�h)��}�(h G@��l߫�h!G��kX�8�Lub�end�h)��}�(h G@\b�-TTh!G��#G�ub�dPivot�h)��}�(h G@\b�-TTh!G��#G�ub�dEnd�h)��}�(h G��Y�+� h!G?�Y�+ˀub�dA�hA)��}�(hDG?Lm��l hEG?Lm���_�hFG?���5�f�ub�dS�G?��N���angleOffset�G��DԂ�length�G@�|��ub�mode�K�active���obj�jj  ub�newObj�h��
startPoint�h)��}�(h G?�uPuPh!G���_�_ubj;  h)��}�(h K h!K ubjP  K �	processed���oldObjectAnchor�h)��}�(h G        h!G        ub�oldObjectAngle�hA)��}�(hDG        hEG        hFG?�      ub�oldObjectScale�G?�      ubj  )��}�(j  j  hj  j   jj  j!  h�ubj  �ComSetBodyAsCurrent���)��}�(j  j  hh�prev�jj  ubj  �ComLoadTexture���)��}�(hj  �newPath�j  �destChannel�K �newSize�j   �oldPath�j  �oldSize�j  ubji  )��}�(hj  jl  j  jm  Kjn  j  jo  j  jp  j  ubj  �ComAddNewShape���)��}�(j  j  hj  �shape�hM�	prevShape�NjN  hubj  �ComNewShapeAddPoint���)��}�(jw  hM�point�hpubjz  )��}�(jw  hMj}  hvubjz  )��}�(jw  hMj}  h|ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubjz  )��}�(jw  hMj}  h�ubj  �ComSelectNextBody���)��}�(j  j  �oldBody�h�oldShape�hM�newBody�h��newShape�N�executed��ubjt  )��}�(j  j  hj  jw  j  jx  NjN  h�ubj�  )��}�(j  j  j�  h�j�  j  j�  jj  j�  Nj�  �ubjt  )��}�(j  j  hj  jw  j�  jx  NjN  jj  ubjd  )��}�(j  j  hh�jg  jj  ubj%  )��}�(h,j+  jS  h�jT  h)��}�(h G?���k���h!G?�HY�^yDubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G        h!G        ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubjd  )��}�(j  j  hjl  jg  h�ubj%  )��}�(h,j+  jS  jj  jT  h)��}�(h G?��KU h!G?�}[1Z� ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G        h!G        ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj%  )��}�(h,j+  jS  jj  jT  h)��}�(h G@��l߫�h!G��kX�8�Lubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G@$��W�h!G���N�1�ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj  �ComAddConstraint���)��}�(hj  j  j  j   j�  j!  Nubj  �ComConstraintSetNewBodyA���)��}�(�entity�j�  j�  hj�  Nubj  �ComConstraintSetNewBodyB���)��}�(j�  j�  j�  h�j�  Nubj  �ComSetAnchorBFromCoords���)��}�(j�  j�  �	newXValue�G�T:'0� �	newYValue�G?��]�1	 �	oldXValue�G        �	oldYValue�G        ubj  �ComSetGrooveAFromCoords���)��}�(j�  j�  j�  G��W��[Lj�  G��W�$@j�  G        j�  G        ubj  �ComSetGrooveBFromCoords���)��}�(j�  j�  j�  G��g}�j�  G?��2�j�  G        j�  G        ubj�  )��}�(hj  j  j  j   j�  j!  j�  ubj  �ComSetConstraintAsCurrent���)��}�(j  j  hj�  jg  j�  ubj�  )��}�(j�  j�  j�  hj�  Nubj�  )��}�(j�  j�  j�  h�j�  Nubj�  )��}�(j�  j�  j�  jj  j�  h�ubj�  )��}�(j�  j�  j�  G@���Mj�  G��6��>�4j�  G        j�  G        ubj�  )��}�(j�  j�  j�  G@���Mj�  G?�XpF�I�j�  G        j�  G        ubj�  )��}�(j�  j�  j�  G@	z:�!Pj�  G?�rCaɐj�  G@���Mj�  G?�XpF�I�ubj�  )��}�(j  j  hj�  jg  j�  ubj�  )��}�(j�  j�  j�  G��W��[Lj�  G?�J�y��j�  G��g}�j�  G?��2�ubj�  )��}�(j  j  )��}�(j  jj  j  j�  j  j�  j  Nj  K hh)��}�(hhj�  j�  j�  j�  jE  jF  ububhj�  jg  Nubj�  )��}�(j  j  )��}�(j  h�j  j  j  j�  j  Nj  K hh)��}�(hhj�  j�  j�  j�  jE  jF  ububhj�  jg  Nubj  �ComSetAnchorB���)��}�(j�  j�  j�  G        j�  G        j�  G�T:'0� j�  G?��]�1	 ubj�  )��}�(j  j  hj�  jg  j�  ubj%  )��}�(h,j*  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G����:>Nh!G��ݯ��ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj5  j8  )��}�(j;  h)��}�(h K h!K ubj>  h)��}�(h G�������h!G��!a�p� ubjA  h)��}�(h G��uL"��xh!G?�׏!snpubjD  h)��}�(h G��uL"��xh!G?�׏!snpubjG  h)��}�(h G?�D@��h!G?���gͼubjJ  hA)��}�(hDG���MN�hEG����{X��hFG?�B����ubjM  G?���l�WjN  G�LGw�/'jO  G?�(����vubjP  KjQ  �jR  h�ubjS  jj  jT  h)��}�(h G@pb�3�Rh!G��%��ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G@      h!G��}���zubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubjd  )��}�(j  j  hh�jg  jj  ubj%  )��}�(h,j  jS  h�jT  h)��}�(h G�������h!G��!a�p� ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G����:>Nh!G��ݯ��ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj%  )��}�(h,j*  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G���3��h!G?�0'\��ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj5  j8  )��}�(j;  h)��}�(h K h!K ubj>  h)��}�(h G����co�(h!G?�(���̈ubjA  h)��}�(h G������rLh!G�ݡ���m�ubjD  h)��}�(h G������rLh!G�ݡ���m�ubjG  h)��}�(h G��=H%~�h!G���^t,tubjJ  hA)��}�(hDG?�+'��0hEG?��_��hFG?� [�ubjM  G@��CO�jN  G@� w��jO  G?�UR��'�ubjP  KjQ  �jR  h�ubjS  jj  jT  h)��}�(h G@6�$
=Th!G���' ��ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G@/tN��h!G��	`��ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubjd  )��}�(j  j  )��}�(j  h�j  j  j  Nj  Nj  K hh)��}�(hhj�  j�  j�  j�  jE  jF  ububhh�jg  jj  ubj%  )��}�(h,j<  jS  h�jT  h)��}�(h G����co�(h!G?�(���̈ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G���3��h!G?�0'\��ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj  )��}�(j  j  )��}�(j  h	�
BodyStatic���)��}�(h�Bottom�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G��r)N���h!G��%�`NGububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@6q�F��h!G?�K����Hubububh,h.)��}�(h1h3)��}�(h6G@��:JMh7G?��}qch8G@ �r���h9G���}qch:G@��:JMh;G?�@�dT ubh<h)��}�(h G@ �r���h!G?�@�dT ubh?hA)��}�(hDG��x[� hEG��T��hFG?��o^�H�ubhGG@�.���ubhH]�hf�Static�h�h�BodyStaticPhysics���)��}�(h�h�)��}�(h�h)��}�(h G        h!G        ubh�h)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubh׉ubh�G?�      h�h�)��}�(h�G?�      h�G        h"G        h׉ubh�h�)��}�(h�G?�      h�G        h"G        h׉ubh�h�)��}�(h�G?�      h�G        h"G        h׉ubububj  hJ�Line���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��q�B�`h!G��""$�ڒububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@� H_:fh!G?�+�(���ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hf�Line�hhhi�LineSpec���)��}�(hn]�(h)��}�(hh)��}�(h G����#h!G���J�hubh"h)��}�(h G����#h!G���J�hububh)��}�(hh)��}�(h G��b�C��h!G���Z�}�ubh"h)��}�(h G��b�C��h!G���Z�}�ububh)��}�(hh)��}�(h G����T^�h!G��Tt�3VLubh"h)��}�(h G����T^�h!G��Tt�3VLububh)��}�(hh)��}�(h G?��l�q�h!G�����/�ubh"h)��}�(h G?��l�q�h!G�����/�ububh)��}�(hh)��}�(h G@\�tLh!G��%��[�ubh"h)��}�(h G@\�tLh!G��%��[�ububh)��}�(hh)��}�(h G@�+�<{Zh!G����Dװubh"h)��}�(h G@�+�<{Zh!G����Dװububh)��}�(hh)��}�(h G@�:GrK�h!G���v�3�ubh"h)��}�(h G@�:GrK�h!G���v�3�ububh)��}�(hh)��}�(h G@8p��h!G��iq�4ubh"h)��}�(h G@8p��h!G��iq�4ububh)��}�(hh)��}�(h G@�|���>h!G���e�.�@ubh"h)��}�(h G@�|���>h!G���e�.�@ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�hŌLinePhysics���)��}�(h�h�)��}�(h�h)��}�(h G?�Ѯ�h!G��Z�5�zubh�h)��}�(h G        h!G        ubh"h)��}�(h G?�Ѯ�h!G��Z�5�zubh׉ubh�G?�S�����h�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G?�      h�G        h"G?�S�����h׉ubh�h�)��}�(h�G?��5^���h�G        h"G?��5^���h׉ubububj  j�  j  j�  j  Khh)��}�(hhj�  j�  j�  j�  jE  jF  ububhj
  j   jr  j!  jj  ubjd  )��}�(j  jn  h�WHeelR_1�jg  jr  ubjd  )��}�(j  jn  hj  jg  jr  ubjd  )��}�(j  jn  hj  jg  jr  ubj%  )��}�(h,j*  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G���qSh!G�Xl"p�pubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj5  j8  )��}�(j;  h)��}�(h K h!K ubj>  h)��}�(h G�X2h!G�=g���ubjA  h)��}�(h G���o�lh!G���<���ubjD  h)��}�(h G���o�lh!G���<���ubjG  h)��}�(h G?���ڀ�4h!G?�fi"$ubjJ  hA)��}�(hDG?��^�X@hEG?�����EhFG?�:	�2xubjM  G?� �����jN  G�O+��jO  G@ȱ�5�ubjP  KjQ  �jR  jr  ubjS  jr  jT  h)��}�(h G@(]��1�Uh!G?�O����,ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G        h!G        ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj  �ComRenameBody���)��}�(jN  jr  hj
  �newName�jt  �oldName�j  ubjt  )��}�(j  jn  hj
  jw  j�  jx  NjN  jr  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubj%  )��}�(h,j  jS  jr  jT  h)��}�(h G�X2h!G�=g���ubj;  h)��}�(h K h!K ubjP  KjY  �jZ  h)��}�(h G���qSh!G�Xl"p�pubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj�  )��}�(j  j  )��}�(j  jr  j  j�  j  j2  j  j�  j  Khh)��}�(hhj�  j�  j�  j�  jE  jF  ububhj�  jg  j�  ubj�  )��}�(hj]  j  j[  j   j�  �DampedRotarySpring���)��}�(h�	CNSTRNT_2�hf�Rotary Spring�j�  Nj�  Nj�  �j�  G?�      �	restAngle�h�UnboundAngle���)��}�(hDG        hEG        hFG?�      ubj  G?�      j   G?�      ubj!  j�  ubj�  )��}�(hj]  j  j[  j   jb  )��}�(h�	CNSTRNT_3�hfjf  j�  Nj�  Nj�  �j�  G?�      jg  ji  )��}�(hDG        hEG        hFG?�      ubj  G?�      j   G?�      ubj!  jc  ubj  �ComDelConstraint���)��}�(hj]  j  j[  j   jn  �objIndex�Kubjt  )��}�(hj]  j  j[  j   jc  jw  Kubj�  )��}�(hj]  j  j[  j   j  j!  j�  ubj�  )��}�(hj]  j  j[  j   j2  j!  j  ubj�  )��}�(j  j[  hj  jg  j2  ubj�  )��}�(j�  j  j�  hj�  Nubj�  )��}�(j�  j  j�  h�j�  Nubj  �ComSetAnchorAFromCoords���)��}�(j�  j  j�  G��W���j�  G���X��j�  G        j�  G        ubj�  )��}�(j�  j  j�  G���A۶j�  G?�����j�  G��W���j�  G���X��ubj�  )��}�(j�  j  j�  G���A۶j�  G?�����j�  G���A۶j�  G?�����ubj�  )��}�(j�  j  j�  G���l�QRj�  G?�dN�f�j�  G���A۶j�  G?�����ubj�  )��}�(j�  j  j�  G���A۶j�  G?䯱��j�  G���l�QRj�  G?�dN�f�ubj�  )��}�(j�  j  j�  G�����Jj�  G?���8߬Hj�  G���A۶j�  G?䯱��ubj�  )��}�(j�  j  j�  G��dn} �j�  G?䯱��j�  G�����Jj�  G?���8߬Hubj�  )��}�(j�  j  j�  G���Àj�  G?䯱��j�  G��dn} �j�  G?䯱��ubj�  )��}�(j�  j  j�  G�:��~b�j�  G����|�xj�  G���Àj�  G?䯱��ubj�  )��}�(j�  j  j�  G���Àj�  G?�����j�  G�:��~b�j�  G����|�xubj�  )��}�(j�  j  j�  G���Àj�  G?�����j�  G���Àj�  G?�����ubj  �ComSetRestLengthFromCoords���)��}�(�newValue�G?����*�j�  j  �oldValue�G?�      ubj�  )��}�(j�  G?���D&�j�  j  j�  G?����*�ubj�  )��}�(j�  G?�/a��Y�j�  j  j�  G?���D&�ubj�  )��}�(j�  G?�� �F j�  j  j�  G?�/a��Y�ubj  �ComSetRestLength���)��}�(j�  j  j�  G        j�  G?�� �F ubj�  )��}�(j  j[  hj4  jg  j  ubj�  )��}�(j�  j2  j�  hj�  Nubj�  )��}�(j�  j2  j�  h�j�  Nubj�  )��}�(j�  j2  j�  jj  j�  h�ubj�  )��}�(j�  j2  j�  G@�[�e�j�  G?�����j�  G        j�  G        ubj�  )��}�(j�  j2  j�  G@�[�e�j�  G?�����M�j�  G@�[�e�j�  G?�����ubj�  )��}�(j�  j2  j�  G@�[�e�j�  G?�����M�j�  G@�[�e�j�  G?�����M�ubj�  )��}�(j�  j2  j�  G        j�  G?�      ubjd  )��}�(j  j  )��}�(j  jr  j  j�  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G��r)N���h!G��%�`NGububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@6q�F��h!G?�K����Hubububh,h.)��}�(h1h3)��}�(h6G@��:JMh7G?��}qch8G@ �r���h9G���}qch:G@��:JMh;G?�@�dT ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hf�Line�hhj�  )��}�(hn]�(h)��}�(hh)��}�(h G�&掷��h!G���/g��Hubh"h)��}�(h G�6YV�4Eh!G���	3^ububh)��}�(hh)��}�(h G@!� �NRh!G� �*-\ubh"h)��}�(h G@5ۍg���h!G��N�[��ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�j�  )��}�(h�h�)��}�(h�h)��}�(h G��{�jb�h!G������ ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��{�jb�h!G������ ubh׉ubh�G?٤��Z1Dh�h�)��}�(h�G?�      h�G        h"G?�      h׉ubh�h�)��}�(h�G?�      h�G        h"G?٤��Z1Dh׉ubh�h�)��}�(h�G@*��՚$�h�G        h"G@*��՚$�h׉ubububj  j2  j  j�  j  Khh)��}�(hhj�  j�  j�  j�  jE  jF  ububhjt  jg  jr  ubj  �ComDelNewShape���)��}�(hj�  j  j�  hj�  jw  j�  �parent�jr  ubjt  )��}�(j  j�  hj�  jw  j�  jx  j�  jN  jr  ubjz  )��}�(jw  j�  j}  j�  ubjz  )��}�(jw  j�  j}  j�  ubj  �ComSetPivot���)��}�(j;  h)��}�(h G?���9~� h!G��<xSm�ub�newWorld�h)��}�(h G?���9~� h!G��<xSm�ub�oldWorld�h)��}�(h K h!K ububj%  )��}�(h,j*  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G@ 5S���&h!G?�	�Ґubh?hA)��}�(hDG        hEG        hFG?�      ubhGG@�.���ubj5  j8  )��}�(j;  h)��}�(h G?���9~� h!G��<xSm�ubj>  h)��}�(h G@9���dc�h!G?��.��E�ubjA  h)��}�(h G@9�0"�jh!G?��X����ubjD  h)��}�(h G@9�<���h!G@Ҝv�ubjG  h)��}�(h G?ґ��� h!G��?Wњc@ubjJ  hA)��}�(hDG��x[� hEG��T��hFG?��o^�H�ubjM  G?�#�`��jN  G?�P��[�jO  G@:G��1�ubjP  K jQ  �jR  jr  ubjS  jr  jT  h)��}�(h G@%�-38�h!G����s=:�ubj;  h)��}�(h G?���9~� h!G��<xSm�ubjP  KjY  �jZ  h)��}�(h G����%<�h!G� ����nubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G?�      ubj%  )��}�(h,j  jS  jr  jT  h)��}�(h G?ɋ9�뎀h!G�#���`ubj;  h)��}�(h G?���9~� h!G��<xSm�ubjP  KjY  �jZ  h)��}�(h G��5�&�jh!G?�	`$��ubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G@�.���ubj%  )��}�(h,j  jS  jr  jT  h)��}�(h G@9���dc�h!G?��.��E�ubj;  h)��}�(h G?���9~� h!G��<xSm�ubjP  K jY  �jZ  h)��}�(h G@ 5S���&h!G?�	�Ґubj]  hA)��}�(hDG        hEG        hFG?�      ubj`  G@�.���ubj�  )��}�(j�  j2  j�  G@=� j�  G��d첾\j�  G@�[�e�j�  G?�����M�ubj�  )��}�(j  j  )��}�(j  jr  j  j�  j  j  j  j�  j  Khh)��}�(hhj�  j�  j�  j�  jE  jF  ububhj  jg  j2  ubj�  )��}�(j�  j  j�  G��i�8j�  G�}��j�  G���Àj�  G?�����ubjd  )��}�(j  j  )��}�(j  jj  j  j�  j  j2  j  j�  j  Khh)��}�(hhj�  j�  j�  j�  jE  jF  ububhjt  jg  jr  ubj  �
ComDelBody���)��}�(hjX  j  jV  j   jr  jw  K�deletedShapes�]�j�  a�constraintsOfDeletedBody�]�ubj  �ComSetStiffness���)��}�(j�  j2  j�  G@@     j�  G?�      ubj  �ComSetDamping���)��}�(j�  j2  j�  G@4      j�  G?�      ubj�  )��}�(j  j  )��}�(j  jj  j  j�  j  j  j  j�  j  Khhubhj  jg  j2  ubjc  )��}�(j�  j  j�  G@@     j�  G?�      ubjg  )��}�(j�  j  j�  G@4      j�  G?�      ubj	  )��}�(j;  h)��}�(h G��t?�լ h!G?�U�ٺ� ubj  h)��}�(h G?]�l%�  h!G�y���D ubj  h)��}�(h K h!K ububj	  )��}�(j;  jt  j  h)��}�(h G?����!�h!G���z�;�ubj  h)��}�(h G?]�l%�  h!G�y���D ububj	  )��}�(j;  jt  j  h)��}�(h G?�l�T��h!G?�����ɀubj  h)��}�(h G?����!�h!G���z�;�ububj	  )��}�(j;  jt  j  h)��}�(h G��t?�լ h!G?�U�ٺ� ubj  h)��}�(h G?�l�T��h!G?�����ɀubube�version��0.0.1�u.