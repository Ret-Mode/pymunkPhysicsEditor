���Z      }�(�database��editorCode.database��Database���)��}�(�bodies�]�(�$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��BODY��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G?u�_�^ h!G?�m��m��ubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�:��:h!G?�PuPuububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]�(�%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?u�_�^ h!G?�������ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�:��:h!G?��m��m�ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��
elasticity�G        �friction�G?�      �isSensor���shapeFilterGroup�K �shapeFilterCategory������ �shapeFilterMask������ �type��Polygon��internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G�A�A�h!G?�333330ubh"h)��}�(h G�A�A�h!G?�333330ububh)��}�(hh)��}�(h G@�+�,h!G?�����ubh"h)��}�(h G@�+�,h!G?�����ububh)��}�(hh)��}�(h G@PuPth!G?�333330ubh"h)��}�(h G@PuPth!G?�333330ububh)��}�(hh)��}�(h G@����h!G?��_�Xubh"h)��}�(h G@����h!G?��_�Xububh)��}�(hh)��}�(h G�������h!G?�I$�I$�ubh"h)��}�(h G�������h!G?�I$�I$�ububh)��}�(hh)��}�(h G��+�,h!G?�I$�I$�ubh"h)��}�(h G��+�,h!G?�I$�I$�ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G��k��k{h!G?ֻ"�B�Nub�user�h)��}�(h G        h!G        ubh"h)��}�(h G��k��k{h!G?ֻ"�B�Nub�userDefined��ub�area�G?�����یdensity�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h��ub�mass�h�)��}�(h�G?�      h�G        h"G?������h��ub�moment�h�)��}�(h�G@m.)O	%h�G        h"G@m.)O	%h��ubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��A�@h!G?�������ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�������h!G?�:��:��ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1�hfG        hgG?�      hh�hiK hj����� hk����� hlhmhnhq)��}�(ht]�(h)��}�(hh)��}�(h G��+�+��h!G?�:��:�ubh"h)��}�(h G��+�+��h!G?�:��:�ububh)��}�(hh)��}�(h G���_�_h!G?�:��:�ubh"h)��}�(h G���_�_h!G?�:��:�ububh)��}�(hh)��}�(h G���m��m�h!G?������ubh"h)��}�(h G���m��m�h!G?������ububh)��}�(hh)��}�(h G?쯊����h!G?�_�_�ubh"h)��}�(h G?쯊����h!G?�_�_�ububh)��}�(hh)��}�(h G?�      h!G?�������ubh"h)��}�(h G?�      h!G?�������ububh)��}�(hh)��}�(h G?�      h!G?��m��m�ubh"h)��}�(h G?�      h!G?��m��m�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G?��8�O�+h!G?�x��7��ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?��8�O�+h!G?�x��7��ubh��ubh�G?��Փ�h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G?��Փ�h��ubh�h�)��}�(h�G?���cB�Dh�G        h"G?���cB�Dh��ubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@ PuPuh!G?㙙����ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��+�,h!G?�PuP�ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfG        hgG?�      hh�hiK hj����� hk����� hlhmhnhq)��}�(ht]�(h)��}�(hh)��}�(h G?�������h!G?�������ubh"h)��}�(h G?�������h!G?�������ububh)��}�(hh)��}�(h G?�fffffdh!G?�:��:��ubh"h)��}�(h G?�fffffdh!G?�:��:��ububh)��}�(hh)��}�(h G@:��:��h!G?�A�A�ubh"h)��}�(h G@:��:��h!G?�A�A�ububh)��}�(hh)��}�(h G@I$�I$�h!G?�������ubh"h)��}�(h G@I$�I$�h!G?�������ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G?�8�fM?h!G?��B�?)ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?�8�fM?h!G?��B�?)ubh��ubh�G?�<���bh�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G?�<���bh��ubh�h�)��}�(h�G?�`����6h�G        h"G?�`����6h��ubububehl�Dynamic�h��+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G?����'�h!G?�%��˨ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?����'�h!G?�%��˨ubh��ubh�G@
fgg\Ph�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@
fgg\Ph�G@Y      h"G@Y      h��ubh�h�)��}�(h�G@L���h�G        h"G@L���h��ubububh)��}�(h�BODY_1�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���J��h!G���-w+ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G���J��h9G        h:G?�      h;G���-w+ubh<h)��}�(h G���J��h!G���-w+ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�hJ�Circle���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���J��h!G���-w+ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G���J��h9G        h:G?�      h;G���-w+ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hfG        hgG?�      hh�hiK hj����� hk����� hl�Circle�hnho�
CircleSpec���)��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj�  �radiusVector�h)��}�(h G        h!G        ubh�h�CircleRadius���)��}�(h"G?�      �base�G?�      ub�	drawLines�K ubh�h��CirclePhysics���)��}�(h�h�)��}�(h�h)��}�(h G���J��h!G���-w+ubh�h)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@4      h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubububahljX  h�j[  )��}�(h�h�)��}�(h�h)��}�(h G���J��h!G���-w+ubh�h)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubh��ubh�G@	!�TD-h�h�)��}�(h�G@v��<:�h�G        h"G        h��ubh�h�)��}�(h�G@4      h�G        h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubububh)��}�(h�BODY_2�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��0�K�h!G��$��,ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G?��0�K�h9G        h:G?�      h;G��$��,ubh<h)��}�(h G?��0�K�h!G��$��,ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�j�  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��0�K�h!G��$��,ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G?��0�K�h9G        h:G?�      h;G��$��,ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_4�hfG        hgG?�      hh�hiK hj����� hk����� hlj�  hnj�  )��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj  j�  h)��}�(h G        h!G        ubh�j�  )��}�(h"G?�      j�  G?�      ubj�  K ubh�j�  )��}�(h�h�)��}�(h�h)��}�(h G?��0�K�h!G��$��,ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@4      h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubububahljX  h�j[  )��}�(h�h�)��}�(h�h)��}�(h G?��0�K�h!G��$��,ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubh��ubh�G@	!�TD-h�h�)��}�(h�G@v��<:�h�G        h"G        h��ubh�h�)��}�(h�G@4      h�G        h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ububube�	shapeList�]�(hMh�j  j�  j�  e�constraints�]�(�/editorCode.constraintInternals.editorConstraint��GrooveJoint���)��}�(h�CNSTRNT�hl�Groove��bodyA�h�bodyB�jl  �selfCollide���maxForce�G�      �maxBias�G�      �	errorBias�G?]q5�NZ�grooveA�h�OffsetPoint���)��}�(�offset�h)��}�(h G���A��h!G��}Nc.M�ubhh)��}�(h G���A��h!G��}Nc.M�ubh"h)��}�(h G���휁h!G�������ubub�grooveB�jW  )��}�(jZ  h)��}�(h G���A��h!G���n�;Yubhh)��}�(h G���A��h!G���n�;Yubh"h)��}�(h G���휁h!G?�?�|�ubub�anchorB�jW  )��}�(jZ  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububjJ  )��}�(h�	CNSTRNT_1�hljN  jO  hjP  j�  jQ  �jR  G�      jS  G�      jT  G?]q5�NZjU  jW  )��}�(jZ  h)��}�(h G?���h�h!G�����0��ubhh)��}�(h G?���h�h!G�����0��ubh"h)��}�(h G?�f�v���h!G��!��Qububja  jW  )��}�(jZ  h)��}�(h G?���/�rh!G��2
�:�ubhh)��}�(h G?���/�rh!G��2
�:�ubh"h)��}�(h G?��8J��dh!G?�2m"�@ububjj  jW  )��}�(jZ  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubububjH  �DampedSpring���)��}�(h�	CNSTRNT_2�hl�Damped Spring�jO  hjP  jl  jQ  �jR  G�      jS  G�      jT  G?������͌
restLength�G        �	stiffness�G@È     �damping�G@Y      �anchorA�jW  )��}�(jZ  h)��}�(h G��y?@<~h!G���\�U�ubhh)��}�(h G��y?@<~h!G���\�U�ubh"h)��}�(h G�����T
h!G��fx�|�ububjj  jW  )��}�(jZ  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububj�  )��}�(h�	CNSTRNT_4�hl�Damped Spring�jO  hjP  jl  jQ  �jR  G�      jS  G�      jT  G?�������j�  G        j�  G@È     j�  G@Y      j�  jW  )��}�(jZ  h)��}�(h G��y?@<~h!G���\�U�ubhh)��}�(h G��y?@<~h!G���\�U�ubh"h)��}�(h G�����T
h!G��fx�|�ububjj  jW  )��}�(jZ  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububj�  )��}�(h�	CNSTRNT_3�hlj�  jO  hjP  j�  jQ  �jR  G�      jS  G�      jT  G?�������j�  G        j�  G@È     j�  G@Y      j�  jW  )��}�(jZ  h)��}�(h G?���e�h!G��:��Abubhh)��}�(h G?���e�h!G��:��Abubh"h)��}�(h G?���,8yh!G��ސێububjj  jW  )��}�(jZ  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubububj�  )��}�(h�	CNSTRNT_5�hlj�  jO  hjP  j�  jQ  �jR  G�      jS  G�      jT  G?�������j�  G        j�  G@È     j�  G@Y      j�  jW  )��}�(jZ  h)��}�(h G?���e�h!G��:��Abubhh)��}�(h G?���e�h!G��:��Abubh"h)��}�(h G?���,8yh!G��ސێububjj  jW  )��}�(jZ  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ububube�mappings�]�(�editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�      h!G��      ubh"h)��}�(h G�      h!G��      ububh)��}�(hh)��}�(h G@      h!G��      ubh"h)��}�(h G@      h!G��      ububh)��}�(hh)��}�(h G�      h!G?�      ubh"h)��}�(h G�      h!G?�      ububh)��}�(hh)��}�(h G@      h!G?�      ubh"h)��}�(h G@      h!G?�      ubube�textureSize�]�(K�K`e�anchor�]�(G@X      G@H      e�mappingSize�]�(K�K`e�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@X      h!G@H      ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububj�  )��}�(h�MAP:1�j�  Kj�  jl  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G���J��h9G        h:G?�      h;G���-w+ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G���v\�Lh!G�vO���ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G��ޕ�r10h!G�vO���ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G���v\�Lh!G��d�k�X ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G��ޕ�r10h!G��d�k�X ububej  ]�(K@K@ej  ]�(G@@      G@@      ej  ]�(K@K@ej  ]�(K K ej  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj"  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububj�  )��}�(h�MAP:1_1�j�  Kj�  j�  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G?��0�K�h9G        h:G?�      h;G��$��,ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?�`2��h!G��r�ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@��L��h!G��r�ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G?�`2��h!G��A''��`ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G@��L��h!G��A''��`ububej  ]�(K@K@ej  ]�(G@@      G@@      ej  ]�(K@K@ej  ]�(K K ej  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj"  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubububeub�textureSizes�]�(K�K`��K@K@��K K ��j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e�texturePaths�]�(�data/textures/truck.png��data/textures/wheel1.png�� �j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�h�currentShape�j  �currentConstraint�j�  �currentMapping�jb  �currentMappingChannel�Khh)��}�(hhjD  jE  jF  jG  j�  j�  ububhj�  �object�h�prevCurrent�Nubj�  )��}�(j�  j�  hj�  j�  jl  j�  hubj�  )��}�(j�  j�  hj�  j�  j�  j�  jl  ubj�  �ComLoadTexture���)��}�(hj�  �newPath�j�  �destChannel�K �newSize�j�  �oldPath�j�  �oldSize�j�  ubj�  )��}�(hj�  j�  j�  j�  Kj�  j�  j�  j�  j�  j�  ubj�  �ComCreateMapping���)��}�(j�  j�  hj�  �mapping�j�  �prevMapping�Nubj�  )��}�(j�  j�  hj�  j�  j)  j�  Nubj�  )��}�(j�  j�  hj�  j�  jb  j�  j)  ubj�  �ComSelectPrevBody���)��}�(j�  j�  �oldBody�j�  �oldShape�N�newBody�jl  �newShape�N�executed��ubj�  )��}�(j�  j�  j�  jl  j�  Nj�  hj�  Nj�  �ubj�  �ComAddNewShape���)��}�(j�  j�  hj�  �shape�hM�	prevShape�Nj�  hubj�  �ComSetNewShapeAsCurrent���)��}�(j�  j�  �newShapeLabel�he�oldShapeLabel�heubj�  �ComNewShapeAddPoint���)��}�(j�  hM�point�hvubj�  )��}�(j�  hMj�  h|ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  j�  hj�  j�  h�j�  hMj�  hubj�  )��}�(j�  j�  j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  j�  hj�  j�  j  j�  h�j�  hubj�  )��}�(j�  j  j�  j.  ubj�  )��}�(j�  j  j�  j4  ubj�  )��}�(j�  j  j�  j:  ubj�  )��}�(j�  j  j�  j@  ubj�  �ComSelectNextBody���)��}�(j�  j�  j�  hj�  j  j�  jl  j�  Nj�  �ubj�  )��}�(j�  j�  hj�  j�  j�  j�  Nj�  jl  ubj�  �ComSetUserParam���)��}�(�param�j�  �oldUserFlag���
oldUserVal�G        �value�G@4      ubj  )��}�(j�  j�  j�  jl  j�  j�  j�  j�  j�  Nj�  �ubj�  )��}�(j�  j�  hj�  j�  j�  j�  Nj�  j�  ubj  )��}�(j"  j0  j#  �j$  G        j%  G@4      ubj�  �ComSetPivot���)��}�(�pivot�h)��}�(h G?��m��h!G��2E\xub�newWorld�h)��}�(h G�����IW~h!G��2E\xub�oldWorld�h)��}�(h K h!K ububj�  �ComSetBodyAsCurrent���)��}�(j�  j�  hjn  �prev�j�  ubj�  �ComStartTransform���)��}�(h,�editorCode.editorViewTransform��ContinuousTransform���)��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�
mouseParam��editorCode.editorMousePivot��MousePivotParams���)��}�(j0  h)��}�(h G?��m��h!G��2E\xub�begin�h)��}�(h G?�Pd?/Fh!G?ޟZؓub�end�h)��}�(h G@��&�Ih!G�������ub�dPivot�h)��}�(h G?�Gu�Gxh!G?���x�8ub�dEnd�h)��}�(h G?��0�K�h!G��$��,ub�dA�hA)��}�(hDG��VlJ�hEG���"(r��hFG��� s�ub�dS�G?�E�����angleOffset�G@ <��P��length�G?�ܪ��<rub�mode�K�active���obj�j�  ub�newObj�jl  �
startPoint�h)��}�(h G?��ư�h!G?�?%�{bDubj0  h)��}�(h G�����IW~h!G��2E\xubji  K�	processed���oldObjectAnchor�h)��}�(h G        h!G        ub�oldObjectAngle�hA)��}�(hDG        hEG        hFG?�      ub�oldObjectScale�G?�      ubj-  )��}�(j0  j1  j3  h)��}�(h G?��m��h!G��2E\xubj6  h)��}�(h G�����IW~h!G��2E\xububj?  )��}�(h,jE  jl  jl  jm  h)��}�(h G?�Ϸ�x�h!G?՗%�<�(ubj0  h)��}�(h G?��m��h!G��2E\xubji  Kjr  �js  h)��}�(h G���J��h!G���-w+ubjv  hA)��}�(hDG        hEG        hFG?�      ubjy  G?�      ubj:  )��}�(j�  j�  hjn  j=  jl  ubj:  )��}�(j�  j�  hj�  j=  jl  ubj?  )��}�(h,jE  jl  j�  jm  h)��}�(h G?�Pd?/Fh!G?ޟZؓubj0  h)��}�(h G?��m��h!G��2E\xubji  Kjr  �js  h)��}�(h G        h!G        ubjv  hA)��}�(hDG        hEG        hFG?�      ubjy  G?�      ubj�  �ComAddConstraint���)��}�(hj�  j�  j�  j�  jK  j�  Nubj�  �ComConstraintSetNewBodyA���)��}�(�entity�jK  j�  hj�  Nubj�  �ComConstraintSetNewBodyB���)��}�(j�  jK  j�  jl  j�  Nubj�  )��}�(j�  jK  j�  j�  j�  jl  ubj�  )��}�(j�  jK  j�  jl  j�  j�  ubj�  �ComSetGrooveAFromCoords���)��}�(j�  jK  �	newXValue�G���A���	newYValue�G��}Nc.M��	oldXValue�G        �	oldYValue�G        ubj�  �ComSetGrooveBFromCoords���)��}�(j�  jK  j�  G���A��j�  G���n�;Yj�  G        j�  G        ubj�  �ComConstraintClone���)��}�(hj�  j�  j�  �baseConstraint�jK  �newConstraint�js  �index�K ubj�  �ComSetConstraintAsCurrent���)��}�(j�  j�  hju  j=  js  ubj�  )��}�(j�  js  j�  j�  j�  jl  ubj�  )��}�(j�  js  j�  G?���/�rj�  G��2
�:�j�  G���A��j�  G���n�;Yubj�  )��}�(j�  js  j�  G?���h�j�  G�����0��j�  G���A��j�  G��}Nc.M�ubj�  )��}�(hj�  j�  j�  j�  j�  j�  js  ubj�  )��}�(j�  j�  j�  hj�  Nubj�  )��}�(j�  j�  j�  jl  j�  Nubj�  �ComSetAnchorAFromCoords���)��}�(j�  j�  j�  G��~���j�  G��kr�uj�  G        j�  G        ubj�  )��}�(j�  j�  j�  G���{6bj�  G��Qk��F�j�  G��~���j�  G��kr�uubj�  )��}�(j�  j�  j�  G��y?@<~j�  G��O�1n�j�  G���{6bj�  G��Qk��F�ubj�  )��}�(j�  j�  j�  G��SJr�j�  G��O�1n�j�  G��y?@<~j�  G��O�1n�ubj�  )��}�(j�  j�  j�  G��SJr�j�  G��O�1n�j�  G��SJr�j�  G��O�1n�ubj�  )��}�(j�  j�  j�  G��ŷ+�Ej�  G��9�He[�j�  G��SJr�j�  G��O�1n�ubj�  )��}�(j�  j�  j�  G���{6bj�  G�� O3:j�  G��ŷ+�Ej�  G��9�He[�ubj�  )��}�(j�  j�  j�  G��y?@<~j�  G���\�U�j�  G���{6bj�  G�� O3:ubj�  �ComSetRestLength���)��}�(j�  j�  �newValue�G        �oldValue�G?�      ubj�  )��}�(hj�  j�  j�  j�  j�  j�  j�  j�  Kubj�  )��}�(j�  j�  j�  j�  j�  jl  ubj�  )��}�(j�  j�  j�  G?���e�j�  G��:��Abj�  G��y?@<~j�  G���\�U�ubj�  �ComSetErrorBias���)��}�(�
constraint�j�  �oldVal�G?]q5�NZ�newVal�G?�������ubj�  �ComSetDamping���)��}�(j�  j�  j�  G@È     j�  G?�      ubj�  �ComSetStiffness���)��}�(j�  j�  j�  G@È     j�  G?�      ubj�  )��}�(j�  j�  hj�  j=  j�  ubj�  )��}�(j�  j�  j�  G@È     j�  G?�      ubj�  )��}�(j�  j�  j�  G@È     j�  G?�      ubj�  )��}�(j�  j�  j�  G?]q5�NZj�  G?�������ubj:  )��}�(j�  j�  hhj=  j�  ubj  )��}�(j"  jh  j#  �j$  G        j%  G@�@     ubj�  )��}�(j�  j�  )��}�(j�  hj�  j  j�  j�  j�  jb  j�  Khhubj�  j  j�  j  ubj�  �ComNewShapeClone���)��}�(hhj�  j  �	baseShape�j�  j�  j�  j�  K j�  j�  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?���D�Ԁh!G��C�S�lububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�������ubububh,h.)��}�(h1h3)��}�(h6G���vf2�hh7G?���6�Ƌh8G?���D�Ԁh9G����6�Ƌh:G���vf2�hh;G��C�S�lubh<h)��}�(h G?���D�Ԁh!G��C�S�lubh?hA)��}�(hDG�c&h�ʐhEG����6�ƋhFG���vf2�hubhGG?�      ubh�SHAPE_5�hfG        hgG?�      hh�hiK hj����� hk����� hlj�  hnj�  )��}�(ht]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G?���D�Ԁh!G��C�S�lububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj*  j�  h)��}�(h G        h!G        ubh�j�  )��}�(h"G?�������j�  G?�      ubj�  K ubh�j�  )��}�(h�h�)��}�(h�h)��}�(h G?���D�Ԁh!G��C�S�lubh�h)��}�(h G        h!G        ubh"h)��}�(h G?���D�Ԁh!G��C�S�lubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@4      h"G@4      h��ubh�h�)��}�(h�G@#������h�G        h"G@#������h��ububububj?  )��}�(h,jD  )��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G��p��
=ph!G?��L��ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubjO  jR  )��}�(j0  h)��}�(h K h!K ubjW  h)��}�(h G?����^�h!G?���m��XubjZ  h)��}�(h G��A��h!G���� �ubj]  h)��}�(h G��A��h!G���� �ubj`  h)��}�(h G���r�8�Th!G��h]5�&Jubjc  hA)��}�(hDG�c&h�ʐhEG����6�ƋhFG���vf2�hubjf  G?�N4�26jg  G?���o�Zjh  G?�d^�ubji  K jj  �jk  j  ubjl  j  jm  h)��}�(h G?���K���h!G?旫Et�bubj0  h)��}�(h K h!K ubji  Kjr  �js  h)��}�(h G        h!G        ubjv  hA)��}�(hDG        hEG        hFG?�      ubjy  G?�      ubj?  )��}�(h,jL  jl  j  jm  h)��}�(h G?����^�h!G?���m��Xubj0  h)��}�(h K h!K ubji  K jr  �js  h)��}�(h G��p��
=ph!G?��L��ubjv  hA)��}�(hDG        hEG        hFG?�      ubjy  G?�      ubj�  �ComDelNewShape���)��}�(hhj�  j  h�SHAPE_5�j�  j  �parent�j�  ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(hhj�  j  j�  j�  j�  j�  j�  Kubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(hhj�  j  j�  j�  j�  j�  j�  Kubj:  )��}�(j�  j  hhj=  j�  ubj  )��}�(j"  jh  j#  �j$  G@�@     j%  G@Y      ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j�  j�  G@Y      j�  G@È     ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j�  j�  G@Y      j�  G@È     ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j�  j�  G@Y      j�  G@È     ubj�  )��}�(j�  j  hj�  j=  j�  ubj�  )��}�(j�  j�  j�  G@Y      j�  G@È     ube�version��0.0.2�u.