��	      }�(�database��editorCode.database��Database���)��}�(�bodies�]��$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��BODY��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G���K�Wk�h!G?�Ƅ��Tubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�Io%�h!G?����l�\ububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?փ��22�r0c1�G��֖�W�r0c2�G��nu�r1c0�G?�֖�W�r1c1�G?փ��22�r1c2�G?ˏ�9�Eub�objectAnchor�h)��}�(h G��nuh!G?ˏ�9�Eub�objectAngle�h�Angle���)��}�(�angle�G?�������sin�G?�Hc�cos�G?����/ub�objectScale�G?��rub�shapes�]��%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���K�Wk�h!G?�Ƅ��Tububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�Io%�h!G?����l�]ubububh,h.)��}�(h1h3)��}�(h6G?փ��22h7G��֖�Wh8G��nuh9G?�֖�Wh:G?փ��22h;G?ˏ�9�Eubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��type��Polygon��internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G��+�+�h!G?ޠ���ubh"h)��}�(h G����#.h!G?��*��OJububh)��}�(hh)��}�(h G?ʃ�:��8h!G?�|W�|W�ubh"h)��}�(h G��Ǟ�L&h!G?�:�L��ububh)��}�(hh)��}�(h G?��A�Bh!G?�PuPtubh"h)��}�(h G���zvLh!G?�[z5���ububh)��}�(hh)��}�(h G?�������h!G?�:��:��ubh"h)��}�(h G��Ԕ֑Eh!G?�[�fububh)��}�(hh)��}�(h G?֠���h!G?�A�A�ubh"h)��}�(h G��,�8�f�h!G?�
wI�ububh)��}�(hh)��}�(h G��������h!G?�A�A� ubh"h)��}�(h G���8�Uqh!G?���L\�6ububh)��}�(hh)��}�(h G������h!G?�uPuPubh"h)��}�(h G�� �8��h!G?�4�sPubube�currentPoint�N�radius�h�Radius���)��}�h"G?�      sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G��ژ?4�h!G?׌m�Sm@ub�user�h)��}�(h G        h!G        ubh"h)��}�(h G��ژ?4�h!G?׌m�Sm@ub�userDefined��ub�area�G@zul�w،density�h�UserSettableFloat���)��}�(h�G?P      h�G        h"G?P      h��ub�mass�h�)��}�(h�G?�      h�G        h"G?szul�w�h��ub�moment�h�)��}�(h�G?"_"wEHh�G        h"G?"_"wEHh��ubububahf�Dynamic�h��+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G��ژ?4�h!G?׌m�Sm@ubh�h)��}�(h G        h!G        ubh"h)��}�(h G��ژ?4�h!G?׌m�Sm@ubh��ubh�G@zul�w�h�h�)��}�(h�G?P      h�G        h"G?P      h��ubh�h�)��}�(h�G?szul�w�h�G        h"G?szul�w�h��ubh�h�)��}�(h�G?"_"wEHh�G        h"G?"_"wEHh��ubububa�	shapeList�]�hMa�constraints�]��mappings�]��editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?փ��22h7G��֖�Wh8G��nuh9G?�֖�Wh:G?փ��22h;G?ˏ�9�Eubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G����_��h!G����Ppd{ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G��{ �:�h!G?�����`ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G��%	�zh!G?��摜�ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G�,1w2h!G?���POiubube�textureSize�]�(K�K`e�anchor�]�(G@X      G@H      e�mappingSize�]�(K*K(e�mappingOffset�]�(KIK,e�uv�]�(h)��}�(h G?�UUUUUUh!G?�UUUUUUubh)��}�(h G?�*�����h!G?�UUUUUUubh)��}�(h G?�UUUUUUh!G?�      ubh)��}�(h G?�*�����h!G?�      ubeh�h)��}�(h G@X�y�E�ah!G@M� ��ub�	subAnchor�h)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G����H�sh!G?�\a�46Jubububaub�textureSizes�]�(K�K`��K K ��j"  j"  j"  j"  j"  j"  j"  j"  j"  j"  j"  j"  j"  j"  e�texturePaths�]�(�data/textures/pinky.png�� �j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  eu.