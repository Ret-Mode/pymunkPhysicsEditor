���K      }�(�database��editorCode.database��Database���)��}�(�bodies�]�(�$editorCode.shapeInternals.editorBody��BodyDynamic���)��}�(�label��BODY��box��editorCode.editorTypes��BoundingBox���)��}�(�center�h�EditorPoint���)��}�(�local�h�V2���)��}�(�x�K �y�K ub�final�h)��}�(h G?u�_�^ h!G?�m��m��ubub�halfWH�h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�:��:h!G?�PuPuububub�	transform�h�ContainerTransform���)��}�(�mat�h�Mat���)��}�(�r0c0�G?�      �r0c1�G�       �r0c2�G        �r1c0�G        �r1c1�G?�      �r1c2�G        ub�objectAnchor�h)��}�(h G        h!G        ub�objectAngle�h�Angle���)��}�(�angle�G        �sin�G        �cos�G?�      ub�objectScale�G?�      ub�shapes�]�(�%editorCode.shapeInternals.editorShape��Polygon���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?u�_�^ h!G?�������ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@�:��:h!G?��m��m�ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE��
elasticity�G        �friction�G?�      �isSensor���shapeFilterGroup�K �shapeFilterCategory������ �shapeFilterMask������ �type�hK�internal��)editorCode.shapeInternals.editorShapeSpec��PolygonSpec���)��}�(�points�]�(h)��}�(hh)��}�(h G�A�A�h!G?�333330ubh"h)��}�(h G�A�A�h!G?�333330ububh)��}�(hh)��}�(h G@�+�,h!G?�����ubh"h)��}�(h G@�+�,h!G?�����ububh)��}�(hh)��}�(h G@PuPth!G?�333330ubh"h)��}�(h G@PuPth!G?�333330ububh)��}�(hh)��}�(h G@����h!G?��_�Xubh"h)��}�(h G@����h!G?��_�Xububh)��}�(hh)��}�(h G�������h!G?�I$�I$�ubh"h)��}�(h G�������h!G?�I$�I$�ububh)��}�(hh)��}�(h G��+�,h!G?�I$�I$�ubh"h)��}�(h G��+�,h!G?�I$�I$�ubube�currentPoint�N�radius�h�Radius���)��}�h"G?�z�G�{sbub�physics��,editorCode.shapeInternals.editorShapePhysics��PolygonPhysics���)��}�(�cog�h�CenterOfGravity���)��}�(�calc�h)��}�(h G��k��k{h!G?ֻ"�B�Nub�user�h)��}�(h G        h!G        ubh"h)��}�(h G��k��k{h!G?ֻ"�B�Nub�userDefined��ub�area�G?�����یdensity�h�UserSettableFloat���)��}�(h�G?�      h�G        h"G?�      h��ub�mass�h�)��}�(h�G?�      h�G        h"G?������h��ub�moment�h�)��}�(h�G@m.)O	%h�G        h"G@m.)O	%h��ubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��A�@h!G?�������ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�������h!G?�:��:��ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_1�hfG        hgG?�      hh�hiK hj����� hk����� hlhKhmhp)��}�(hs]�(h)��}�(hh)��}�(h G��+�+��h!G?�:��:�ubh"h)��}�(h G��+�+��h!G?�:��:�ububh)��}�(hh)��}�(h G���_�_h!G?�:��:�ubh"h)��}�(h G���_�_h!G?�:��:�ububh)��}�(hh)��}�(h G���m��m�h!G?������ubh"h)��}�(h G���m��m�h!G?������ububh)��}�(hh)��}�(h G?쯊����h!G?�_�_�ubh"h)��}�(h G?쯊����h!G?�_�_�ububh)��}�(hh)��}�(h G?�      h!G?�������ubh"h)��}�(h G?�      h!G?�������ububh)��}�(hh)��}�(h G?�      h!G?��m��m�ubh"h)��}�(h G?�      h!G?��m��m�ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G?��8�O�+h!G?�x��7��ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?��8�O�+h!G?�x��7��ubh��ubh�G?��Փ�h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G?��Փ�h��ubh�h�)��}�(h�G?���cB�Dh�G        h"G?���cB�Dh��ubububhL)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G@ PuPuh!G?㙙����ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��+�,h!G?�PuP�ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_2�hfG        hgG?�      hh�hiK hj����� hk����� hlhKhmhp)��}�(hs]�(h)��}�(hh)��}�(h G?�������h!G?�������ubh"h)��}�(h G?�������h!G?�������ububh)��}�(hh)��}�(h G?�fffffdh!G?�:��:��ubh"h)��}�(h G?�fffffdh!G?�:��:��ububh)��}�(hh)��}�(h G@:��:��h!G?�A�A�ubh"h)��}�(h G@:��:��h!G?�A�A�ububh)��}�(hh)��}�(h G@I$�I$�h!G?�������ubh"h)��}�(h G@I$�I$�h!G?�������ububeh�Nh�h�)��}�h"G?�z�G�{sbubh�h�)��}�(h�h�)��}�(h�h)��}�(h G?�8�fM?h!G?��B�?)ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?�8�fM?h!G?��B�?)ubh��ubh�G?�<���bh�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G        h"G?�<���bh��ubh�h�)��}�(h�G?�`����6h�G        h"G?�`����6h��ubububehl�Dynamic�h��+editorCode.shapeInternals.editorBodyPhysics��BodyPhysics���)��}�(h�h�)��}�(h�h)��}�(h G?����'�h!G?�%��˨ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?����'�h!G?�%��˨ubh��ubh�G@
fgg\Ph�h�)��}�(h�G?�      h�G        h"G        h��ubh�h�)��}�(h�G@
fgg\Ph�G@�@     h"G@�@     h��ubh�h�)��}�(h�G@L���h�G        h"G@L���h��ubububh)��}�(h�BODY_1�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���J��h!G���-w+ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G���J��h9G        h:G?�      h;G���-w+ubh<h)��}�(h G���J��h!G���-w+ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�hJ�Circle���)��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G���J��h!G���-w+ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G���J��h9G        h:G?�      h;G���-w+ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_3�hfG        hgG?�      hh�hiK hj����� hk����� hlj�  hmhn�
CircleSpec���)��}�(hs]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj�  �radiusVector�h)��}�(h G        h!G        ubh�h�CircleRadius���)��}�(h"G?�      �base�G?�      ub�	drawLines�K ubh�h��CirclePhysics���)��}�(h�h�)��}�(h�h)��}�(h G���J��h!G���-w+ubh�h)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@4      h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubububahljW  h�jZ  )��}�(h�h�)��}�(h�h)��}�(h G���J��h!G���-w+ubh�h)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubh��ubh�G@	!�TD-h�h�)��}�(h�G@v��<:�h�G        h"G        h��ubh�h�)��}�(h�G@4      h�G        h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubububh)��}�(h�BODY_2�hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��0�K�h!G��$��,ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G?��0�K�h9G        h:G?�      h;G��$��,ubh<h)��}�(h G?��0�K�h!G��$��,ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubhH]�j�  )��}�(hh)��}�(hh)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?��0�K�h!G��$��,ububh%h)��}�(hh)��}�(h K h!K ubh"h)��}�(h G?�      h!G?�      ubububh,h.)��}�(h1h3)��}�(h6G?�      h7G�       h8G?��0�K�h9G        h:G?�      h;G��$��,ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubh�SHAPE_4�hfG        hgG?�      hh�hiK hj����� hk����� hlj�  hmj�  )��}�(hs]�(h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ububh)��}�(hh)��}�(h G?�      h!G        ubh"h)��}�(h G        h!G        ububehj  j�  h)��}�(h G        h!G        ubh�j�  )��}�(h"G?�      j�  G?�      ubj�  K ubh�j�  )��}�(h�h�)��}�(h�h)��}�(h G?��0�K�h!G��$��,ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubh��ubh�G@	!�TD-h�h�)��}�(h�G?�      h�G        h"G?�      h��ubh�h�)��}�(h�G?�      h�G@4      h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ubububahljW  h�jZ  )��}�(h�h�)��}�(h�h)��}�(h G?��0�K�h!G��$��,ubh�h)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubh��ubh�G@	!�TD-h�h�)��}�(h�G@v��<:�h�G        h"G        h��ubh�h�)��}�(h�G@4      h�G        h"G@4      h��ubh�h�)��}�(h�G@$      h�G        h"G@$      h��ububube�	shapeList�]�(hMh�j  j�  j�  e�constraints�]�(�/editorCode.constraintInternals.editorConstraint��GrooveJoint���)��}�(h�CNSTRNT�hl�Groove��bodyA�h�bodyB�jk  �selfCollide���maxForce�G�      �maxBias�G�      �	errorBias�G?]q5�NZ�grooveA�h�OffsetPoint���)��}�(�offset�h)��}�(h G���A��h!G��}Nc.M�ubhh)��}�(h G���A��h!G��}Nc.M�ubh"h)��}�(h G���휁h!G�������ubub�grooveB�jU  )��}�(jX  h)��}�(h G���A��h!G���n�;Yubhh)��}�(h G���A��h!G���n�;Yubh"h)��}�(h G���휁h!G?�?�|�ubub�anchorB�jU  )��}�(jX  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububjH  )��}�(h�	CNSTRNT_1�hljL  jM  hjN  j�  jO  �jP  G�      jQ  G�      jR  G?]q5�NZjS  jU  )��}�(jX  h)��}�(h G?���h�h!G�����0��ubhh)��}�(h G?���h�h!G�����0��ubh"h)��}�(h G?�f�v���h!G��!��Qububj_  jU  )��}�(jX  h)��}�(h G?���/�rh!G��2
�:�ubhh)��}�(h G?���/�rh!G��2
�:�ubh"h)��}�(h G?��8J��dh!G?�2m"�@ububjh  jU  )��}�(jX  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubububjF  �DampedSpring���)��}�(h�	CNSTRNT_2�hl�Damped Spring�jM  hjN  jk  jO  �jP  G�      jQ  G�      jR  G?������͌
restLength�G        �	stiffness�G@È     �damping�G@È     �anchorA�jU  )��}�(jX  h)��}�(h G��y?@<~h!G���\�U�ubhh)��}�(h G��y?@<~h!G���\�U�ubh"h)��}�(h G�����T
h!G��fx�|�ububjh  jU  )��}�(jX  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububj�  )��}�(h�	CNSTRNT_3�hlj�  jM  hjN  j�  jO  �jP  G�      jQ  G�      jR  G?�������j�  G        j�  G@È     j�  G@È     j�  jU  )��}�(jX  h)��}�(h G?���e�h!G��:��Abubhh)��}�(h G?���e�h!G��:��Abubh"h)��}�(h G?���,8yh!G��ސێububjh  jU  )��}�(jX  h)��}�(h G        h!G        ubhh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ububube�mappings�]�(�editorCode.textureMapping��TextureMapping���)��}�(h�MAP:0��channel�K �body�hh,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�mappingRect�]�(h)��}�(hh)��}�(h G�      h!G��      ubh"h)��}�(h G�      h!G��      ububh)��}�(hh)��}�(h G@      h!G��      ubh"h)��}�(h G@      h!G��      ububh)��}�(hh)��}�(h G�      h!G?�      ubh"h)��}�(h G�      h!G?�      ububh)��}�(hh)��}�(h G@      h!G?�      ubh"h)��}�(h G@      h!G?�      ubube�textureSize�]�(K�K`e�anchor�]�(G@X      G@H      e�mappingSize�]�(K�K`e�mappingOffset�]�(K K e�uv�]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@X      h!G@H      ub�	subAnchor�h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G        h!G        ubububj�  )��}�(h�MAP:1�j�  Kj�  jk  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G���J��h9G        h:G?�      h;G���-w+ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G���v\�Lh!G�vO���ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G��ޕ�r10h!G�vO���ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G���v\�Lh!G��d�k�X ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G��ޕ�r10h!G��d�k�X ububej�  ]�(K@K@ej�  ]�(G@@      G@@      ej�  ]�(K@K@ej�  ]�(K K ej�  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G���J��h!G���-w+ubububj�  )��}�(h�MAP:1_1�j�  Kj�  j�  h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G?��0�K�h9G        h:G?�      h;G��$��,ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ubj�  ]�(h)��}�(hh)��}�(h G��      h!G��      ubh"h)��}�(h G?�`2��h!G��r�ububh)��}�(hh)��}�(h G?�      h!G��      ubh"h)��}�(h G@��L��h!G��r�ububh)��}�(hh)��}�(h G��      h!G?�      ubh"h)��}�(h G?�`2��h!G��A''��`ububh)��}�(hh)��}�(h G?�      h!G?�      ubh"h)��}�(h G@��L��h!G��A''��`ububej�  ]�(K@K@ej�  ]�(G@@      G@@      ej�  ]�(K@K@ej�  ]�(K K ej�  ]�(h)��}�(h G        h!G        ubh)��}�(h G?�      h!G        ubh)��}�(h G        h!G?�      ubh)��}�(h G?�      h!G?�      ubeh�h)��}�(h G@@      h!G@@      ubj�  h)��}�(hh)��}�(h G        h!G        ubh"h)��}�(h G?��0�K�h!G��$��,ubububeub�textureSizes�]�(K�K`��K@K@��K K ��jv  jv  jv  jv  jv  jv  jv  jv  jv  jv  jv  jv  jv  e�texturePaths�]�(�data/textures/truck.png��data/textures/wheel1.png�� �j{  j{  j{  j{  j{  j{  j{  j{  j{  j{  j{  j{  j{  e�queueProcessed��collections��deque���)KȆ�R�(�editorCode.commandExec��
ComAddBody���)��}�(�state��editorCode.editorState��EditorState���)��}�(�currentBody�h�currentShape�j  �currentConstraint�j�  �currentMapping�j9  �currentMappingChannel�Khhubhh�object�h�prevCurrent�Nubj�  )��}�(j�  j�  hhj�  jk  j�  hubj�  )��}�(j�  j�  hhj�  j�  j�  jk  ubj�  �ComLoadTexture���)��}�(hh�newPath�jy  �destChannel�K �newSize�jt  �oldPath�j{  �oldSize�jv  ubj�  )��}�(hhj�  jz  j�  Kj�  ju  j�  j{  j�  jv  ubj�  �ComCreateMapping���)��}�(j�  j�  hh�mapping�j�  �prevMapping�Nubj�  )��}�(j�  j�  hhj�  j   j�  Nubj�  )��}�(j�  j�  hhj�  j9  j�  j   ubj�  �ComSelectPrevBody���)��}�(j�  j�  �oldBody�j�  �oldShape�N�newBody�jk  �newShape�N�executed��ubj�  )��}�(j�  j�  j�  jk  j�  Nj�  hj�  Nj�  �ubj�  �ComAddNewShape���)��}�(j�  j�  hh�shape�hM�	prevShape�Nj�  hubj�  �ComSetNewShapeAsCurrent���)��}�(j�  j�  �newShapeLabel�he�oldShapeLabel�heubj�  �ComNewShapeAddPoint���)��}�(j�  hM�point�huubj�  )��}�(j�  hMj�  h{ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  hMj�  h�ubj�  )��}�(j�  j�  hhj�  h�j�  hMj�  hubj�  )��}�(j�  j�  j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  h�j�  h�ubj�  )��}�(j�  j�  hhj�  j  j�  h�j�  hubj�  )��}�(j�  j  j�  j-  ubj�  )��}�(j�  j  j�  j3  ubj�  )��}�(j�  j  j�  j9  ubj�  )��}�(j�  j  j�  j?  ubj�  �ComSelectNextBody���)��}�(j�  j�  j�  hj�  j  j�  jk  j�  Nj�  �ubj�  )��}�(j�  j�  hhj�  j�  j�  Nj�  jk  ubj�  �ComSetUserParam���)��}�(�param�j�  �oldUserFlag���
oldUserVal�G        �value�G@4      ubj�  )��}�(j�  j�  j�  jk  j�  j�  j�  j�  j�  Nj�  �ubj�  )��}�(j�  j�  hhj�  j�  j�  Nj�  j�  ubj�  )��}�(j�  j.  j�  �j�  G        j�  G@4      ubj�  �ComSetPivot���)��}�(�pivot�h)��}�(h G?��m��h!G��2E\xub�newWorld�h)��}�(h G�����IW~h!G��2E\xub�oldWorld�h)��}�(h K h!K ububj�  �ComSetBodyAsCurrent���)��}�(j�  j�  hjm  �prev�j�  ubj�  �ComStartTransform���)��}�(h,�editorCode.editorViewTransform��ContinuousTransform���)��}�(h,h.)��}�(h1h3)��}�(h6G?�      h7G        h8G        h9G        h:G?�      h;G        ubh<h)��}�(h G        h!G        ubh?hA)��}�(hDG        hEG        hFG?�      ubhGG?�      ub�
mouseParam��editorCode.editorMousePivot��MousePivotParams���)��}�(j  h)��}�(h G?��m��h!G��2E\xub�begin�h)��}�(h G?�Pd?/Fh!G?ޟZؓub�end�h)��}�(h G@��&�Ih!G�������ub�dPivot�h)��}�(h G?�Gu�Gxh!G?���x�8ub�dEnd�h)��}�(h G?��0�K�h!G��$��,ub�dA�hA)��}�(hDG��VlJ�hEG���"(r��hFG��� s�ub�dS�G?�E�����angleOffset�G@ <��P��length�G?�ܪ��<rub�mode�K�active���obj�j�  ub�newObj�jk  �
startPoint�h)��}�(h G?��ư�h!G?�?%�{bDubj  h)��}�(h G�����IW~h!G��2E\xubj>  K�	processed���oldObjectAnchor�h)��}�(h G        h!G        ub�oldObjectAngle�hA)��}�(hDG        hEG        hFG?�      ub�oldObjectScale�G?�      ubj  )��}�(j  j  j  h)��}�(h G?��m��h!G��2E\xubj  h)��}�(h G�����IW~h!G��2E\xububj  )��}�(h,j  jA  jk  jB  h)��}�(h G?�Ϸ�x�h!G?՗%�<�(ubj  h)��}�(h G?��m��h!G��2E\xubj>  KjG  �jH  h)��}�(h G���J��h!G���-w+ubjK  hA)��}�(hDG        hEG        hFG?�      ubjN  G?�      ubj  )��}�(j�  j�  hjm  j  jk  ubj  )��}�(j�  j�  hj�  j  jk  ubj  )��}�(h,j  jA  j�  jB  h)��}�(h G?�Pd?/Fh!G?ޟZؓubj  h)��}�(h G?��m��h!G��2E\xubj>  KjG  �jH  h)��}�(h G        h!G        ubjK  hA)��}�(hDG        hEG        hFG?�      ubjN  G?�      ubj�  �ComAddConstraint���)��}�(hhj�  j�  j�  jI  j�  Nubj�  �ComConstraintSetNewBodyA���)��}�(�entity�jI  j�  hj�  Nubj�  �ComConstraintSetNewBodyB���)��}�(ju  jI  j�  jk  j�  Nubjw  )��}�(ju  jI  j�  j�  j�  jk  ubjw  )��}�(ju  jI  j�  jk  j�  j�  ubj�  �ComSetGrooveAFromCoords���)��}�(ju  jI  �	newXValue�G���A���	newYValue�G��}Nc.M��	oldXValue�G        �	oldYValue�G        ubj�  �ComSetGrooveBFromCoords���)��}�(ju  jI  j�  G���A��j�  G���n�;Yj�  G        j�  G        ubj�  �ComConstraintClone���)��}�(hhj�  j�  �baseConstraint�jI  �newConstraint�jq  �index�K ubj�  �ComSetConstraintAsCurrent���)��}�(j�  j�  hjs  j  jq  ubjw  )��}�(ju  jq  j�  j�  j�  jk  ubj�  )��}�(ju  jq  j�  G?���/�rj�  G��2
�:�j�  G���A��j�  G���n�;Yubj  )��}�(ju  jq  j�  G?���h�j�  G�����0��j�  G���A��j�  G��}Nc.M�ubjn  )��}�(hhj�  j�  j�  j�  j�  jq  ubjr  )��}�(ju  j�  j�  hj�  Nubjw  )��}�(ju  j�  j�  jk  j�  Nubj�  �ComSetAnchorAFromCoords���)��}�(ju  j�  j�  G��~���j�  G��kr�uj�  G        j�  G        ubj�  )��}�(ju  j�  j�  G���{6bj�  G��Qk��F�j�  G��~���j�  G��kr�uubj�  )��}�(ju  j�  j�  G��y?@<~j�  G��O�1n�j�  G���{6bj�  G��Qk��F�ubj�  )��}�(ju  j�  j�  G��SJr�j�  G��O�1n�j�  G��y?@<~j�  G��O�1n�ubj�  )��}�(ju  j�  j�  G��SJr�j�  G��O�1n�j�  G��SJr�j�  G��O�1n�ubj�  )��}�(ju  j�  j�  G��ŷ+�Ej�  G��9�He[�j�  G��SJr�j�  G��O�1n�ubj�  )��}�(ju  j�  j�  G���{6bj�  G�� O3:j�  G��ŷ+�Ej�  G��9�He[�ubj�  )��}�(ju  j�  j�  G��y?@<~j�  G���\�U�j�  G���{6bj�  G�� O3:ubj�  �ComSetRestLength���)��}�(ju  j�  �newValue�G        �oldValue�G?�      ubj�  )��}�(hhj�  j�  j�  j�  j�  j�  j�  Kubjw  )��}�(ju  j�  j�  j�  j�  jk  ubj�  )��}�(ju  j�  j�  G?���e�j�  G��:��Abj�  G��y?@<~j�  G���\�U�ubj�  �ComSetErrorBias���)��}�(�
constraint�j�  �oldVal�G?]q5�NZ�newVal�G?�������ubj�  �ComSetDamping���)��}�(ju  j�  j�  G@È     j�  G?�      ubj�  �ComSetStiffness���)��}�(ju  j�  j�  G@È     j�  G?�      ubj�  )��}�(j�  j�  hj�  j  j�  ubj�  )��}�(ju  j�  j�  G@È     j�  G?�      ubj�  )��}�(ju  j�  j�  G@È     j�  G?�      ubj�  )��}�(j�  j�  j�  G?]q5�NZj�  G?�������ubj  )��}�(j�  j�  hhj  j�  ubj�  )��}�(j�  jg  j�  �j�  G        j�  G@�@     ube�version��0.0.2�u.